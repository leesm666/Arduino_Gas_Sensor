PK   w�X��m  �L    cirkitFile.json�]s�F�����s�[EhЍo�%�Im�6�f+{a�T�b�Mj@ʎ����ݠl��D�}�b=Sq$���y�h6N>κ�]���7]{�����zv����M�5���߆���r}����ڕwof7�����]ԛ�w�u���&m�&UA�ję^U���-�*��&L��6�ݼ|=�\ɚkY�h�y��6-�0(Z]qT�A�(�Iu�y��G���|��Y͇���\�=6Ϳ6�ۼo��+���8L�2�TP�ahZ�UP��H�We�dy��ѭ2��۬�n��`og��$2"��y&k�˚G*T][6��\��J^I�_x(�������텕����2�5~����R^�Υ�R�ҹ\X�ZX�ZX�ZX�ZX�:N���$�K?>}���#a�G��� ���K'��p2�
��m2~��'��K�(vh�i_@�܁desZx��زQl�H�9�l�X��
ѡq�.�J��kVz-\���ř��A������N�N�+����	)~R�ɔ���3���r�c��b�����O��B�H�|�V���O�O���/t���<e�KY����O��B�J�|�3V���O�O���/t���<g��Y����O����S��/X�
V?)?��S,���>f�}�h
���LQ�C�[��N�Z���Z(ES��&G�:�O)ؠST0ES�o�G�:l)�ST0ES���G�:��(ؚST0ES��#F�glЈ)*���)���4
�iz��1?!(T�.!9�;HA�]#�F
�����N;$Tv�������6��},Y�x��囝���6;<���p�b��`+L�
Ȥ i����v��A`'M�N����)*�b�n�1갓�a'MLQ�L1t�F�uz���KL1t7��u�IӰ�&��`�
���	�u�IӰ�&��`�
��/k�u�IӰ�&��`�
���̌u�IӰ�&��`�
��_\�:l_iؾST0ES��	G��4��)*���)��kt#F�}4���)*��z��Wg*��0nE�Qc�6(�Q�(�"��E�?��pV��x�j>��Y���O}{�QoV�N�1�K���y{unB����)�sc; �'��� ��آ|��%A��"(��#(�EI�T�����e�W1嫘�U1�T�bJX�5���oEu��*�Y��b��Lk��5SŚ�b�T��X�\'����j�x!�a�8b�8��Q!> y���/�	�jOڽ��S2�nX�o.�{�hr���
*�v31|�^y�sMܛ�i8*���_'��
�~\��5=�|��Qਠ�u���aT�X���"pTPi��"���J,���8*�4Dڍ��QA����8*�4D���QA�LEyZ�
*�v#,pTP��L�k���JC�ݰTz��'`ਠ�i7G�����aI���	��aI�9�l"�l"��s˦��I܀��3'���%��x{B9xXRo�6sb,xXRo��'���%���3'���%����Ix{�> �1͉��aI�1mޞdHo�Hs�/xXR����MÒzcv��K�Òz���8�����\�L5'F��%�غ�g@zO��25xXR�¿�ˀ���_��	$h���_���']��ל 
����&������6�M�#m�-i��6	oOb�7�9�<,�7�M�ۓ���kNK��k�����@zc����Òzc��$�=y!�ޘ��Dk���^�Ix{�E �1�	��aI��k���d�@zc����Òzc��&��I+����5'؃�%��v�M�ۓk⃽<�@y��s�N �ç���'�]�k��'��~ו+�Ύ>��h%z
���9ʓ�rv���AI�A��A)������^Ŕ�b�W1��
VL	+��SĊ�b�T���`��5SŚ�b�T�f�X3U��*�LGLGU<.��D�Ш�g���H{�OhT����>�QA�!Ҟ�Tz��D�Ш��iO�	�
*=�| �OhTPi��'��F�X��'4*�4D�}B��J,�T"�>�QA�����T"�>�QA�e��T"�>�QA�� ��F��H{�OhTP�C�>�QA�!Ҟ��tN0�̍ �aI���&��>a�欲�����2�-��.��/�J��>�aI�1�l޾�Fo�6s#@pXRo�9���/���3������&��>a��,47�%��\�Ix��O�1#͍ �aI�1/m޾�Fo�Ns#@pXRo�Q���/���3������&��>a�Ƭ57�%��ܵIx��O��*���F����_���/����������&��>a��6�M�#m�-iܞ��6�M��j'�OpXRo�_���/����������&��>a���57�%����Ix��O�1͍ �aI�1m޾�Fo�_s#@pXRo�_���/����������&��>a���57�%����Ix��O<�#�O�(O�5}v���)�������z��t�����M6��_v���nU�ms�\�n���f7/_�>S�i��uTY��J�TiDy['y6Qe?SVy���_���0䘷������Ͽ<"At������+'��QO�h�o��;F`Ot&+[U�>>�(��B��l�P�s��%\ag"Yg�G�r�� ��{iwRvC��ן��]�v�����u�ÿ47'��߂��s��hߞ�c��Vrg)3��z9=�R�|����x?K\ٟE�矏���e�/����t�ϵ�?-�?Y���<��D��OM�O@/�g(y/�R���B�?X!}��^�Y�A�t�~���&�������h��4h��o�1-i�����gJK�?���iI{)�u&<��p��;��}&l���pƒ����>��@��B��'E ҢTҪ�_:)�������Т�iKZ�Z<qJSKSKSKSKS{
SK�r/��I�4��i���l�#��wb8�px�"��$���{�'q!cO��c��Tg�&λ$����'�����`�y8��
�ySD(�vEH0+�pƏuw\t�P�%�8rM�W8�'�G�cg�v�&΋!����'���CTtV˗������(��	^���G��G�y���CTS�*sx����v��;�fpx��b���dQѱ�.u�QQL����!*:���F��!*�)z��9<DE����O�Dn���C���������A�DB,K_4�TK�rcyA@FK1K_�0�h	�=n�.�h)f�-SǍ�-_f��j	X;nT.�h	�;0K_�TK��qcpA@F��5�s��������=[$�=��E�~��#����N�z+U���+#���#�t��	6B	�>r�m��z�e
w�ä}�������ڂ���Q�Y�{�Z��V2Z����+Ւ�V��+�7����+�p�ܐY��p�`��]�����Ȃ��������J�%7d�%��/�V�%�(���  �%�kf���j	xFn�+�h	��Y�Bk�Z���
2Z;�`��@Z���䆱�����>"��/l�pD̬��#�e�-+i���4�}m�ll΁�ڠ�sRf7/g�}.�:���lF����܆�}�;cb�i�>��Ɔ���D{���*{��'+{v�чU(�@�ڶ�=�m�mm[h�B�}2K��m�ȶ����9���mF�~?��vg��֜d�N��~�<�=O���Z��wtf��#:�Ę�_ZHzD$���
z��������z�����ё�������)����҉>_'�J_�U���;�����4�΂�!����{(z8���C�{(y8���҇C�{({8����C�������$��bs�ZnwV���7�/��ww�ު(�>�{�ar�;}{gK�>��T��[��ˋ���^t����-[��1b*d�[n��,�΋4�b�'�Q����0����e�Cc���$4�M�� -�((�E�Q���H�P۴�/����'���,�v�������6�Ҡ����K����U�@�*���`�$�.�į��������������o��ϻ�f��2"3u]G�@="��ޭ�_v�͙�]�\�j��˷�g{t>{W���O���m/���Ҕ��������O����fQ���9�m�_��e�j���k�y��Z#��Ԛ)����~Qֻ��+w�𴃞�#À�Wi%ss}��:9,F5U�Q�%IdqXe�� �"�,��X�U�g-�O��[��f��cT�k��$4=��C\�?d�G��#�����:<�����Ӣ���><����I��:>���0H��q<p@�P-�"w/+�y�Ёt�#�d�E4�B����s ��n/��@2�"j��Z��V��V��+2I�|�Y5m7����z_�n^Ͷ����ͫ���l�����(I���I�?�|��i�$q�FZ�y���o�[m�e�����m����ʃ�����yPfi,�n��m�}[����:�ꬩ�,���YTy�����rm�ŗv?���w��h��UV��4��07����'Յ���������Z�͘��<�|e�ݛ�9@�c�Qk/���U����� YD��T4EZ룡����v}ؿE�	���͂�.��0�:˲2o�EyP�[m��ao��*�&4O�������^�������O<���]�nZ��N��w���U������a���|��ܯ7}����J���t�o��k�ۇc��jnFj�X�ZOq]/�
�)ꅹ͛):Wy/�ʡ��b9,JU�M��l���l��eؚ+�ʂ��lVf�.�67S}ZW���TS�͢��:����R3Amj�l�j�,,0�3��uP���H�ja��QTGU��u�x���_��m��ն����ۿ_}|�j}u�׿^��������G���Woڮ�_�6W���jc�O7�l��O��z��f��y[.����k�]۬>��{�s�j�]_2}�?���l?{��}fxqrN��:;�q�1��㛻�֯sÎ����12u�$1����:Z��uVV��\������ԋ�SdUZ�uzo�����uz�_����/�=�x��>�͡4<��?'K�'׏�Qcs�n�u�nc�Y� SKS�Ӿ��wqqmf���{�lvo��D5��|���s���S���O~8��iY�i�o�<������/������p�}��h�sI���_T^|�mܗ���۽X�.���~�X7,�?�Cw���Ѿ��O�ݻ�r�{Q����f�x5��?-^�?�k�����K�O����sk�k%hϘ�d�Ӳ���/�Ej�iǗ�=��'s+2�y\e���,F���煋,�k���k��8��<�x�NG�ffP�i�S���G+3�U���������b��/��W���ß��q���`tr|��sf�sOK�uu:������6^����OX09]09R0�<��<->o�H�T���nF|��B1]�pD��^^��1��w��g�q��9���b�"������ט��6��Kk.�/ZN���i���#��E�.Z͎�?���t]*r�b�9����G�/�'\kd<�x:/]{8��p�b�@�l	��`>�/O�%��8��� ��[�V?-~,wm�,Wv맩�m���_m�c��/W�n���k�ZO��k[9w���z��v[w˻�r��� PK   w�X�<1	}�  � /   images/02d8db12-ba28-4e49-8e56-db179b980a39.pngԼ�WSY�>�Agl�b�HDz� �H�)�AJBI(c���@��H��B��!TC'�J(��N|�x���keapg�{�庮{�s��=��t^]M�!t�
���)�/�]�ׯ��~~P�Y� ��f�q~��N|�7��x�S屧��SO�'�6 ///a{G�'�l�]�m߭�_���+�5�N^��IN�IY��t�MQ�&���w߻h����wU��p��]���x
o�qOֳUm��C����Iw�M�����_�Fkp�7JQ�:o�V��o�o`��Z��dW#8�Pv�F���*#蟟4��G�cB��ܯ�������?�}���~����;ƺ�N�M�!Pu���%��cS	�=�zl�8�co۟?�;�����\�$�����;|gGo�m�'�ODۏr젩!!�e��H�P3����w�f]����E�k�p{�� �����-7�������� R~	<�����0��,T_�ӑc �r[�k=�[W��uEO�_�]+	}:�պ:zE}=Uo�[�b�5K<�Z�����V�UU�o�zE�<�]f�oQ�.Q�}
�����;�Ue->�\����D]����-��.��I�յ~b�2+��)2�32+wV'�B�kY�@ A��+��⡃A�z�66�L�������;m��ѣ�7�$��]��R�^Q�=�svgn~U�b[��oI�ԉ���x�O��Mr��T߀rR��P�����o񯣼��NbLMYߍ����+�u��G��5�I,�;՚I[�]˯��zXӋ�M*}z���������C��H*s��J�ҳ�k9{%(+��c���_�xu�K�@>iY�����وG��AF���L�Oo�f�q+�T�y<7iX��֣	�6\���o�`Q�F
̆��p�a(c|+|�{َVG�����2����a'�g	p�-��+��=�D��V��(AGN��d<N�#1�v���s-��u)_���	���`"�
��qj7�'4��m[a�,ӰQ�n�<G�ؕ�_�nLI�
��LB��fM��0�W�]ܺ2�H�i[�cSg_p�k8������^���^ٝ�V��L0#H��^>V�GQB����s:�ɺ"=��PV�Nv7q�\�pEE���
%)��f���}�_��~����	K�s;xz]�V�3R��E�`I�@▝ܬ�P����4��uXKV��.�>��4}��S���;�z@�ަ6���ҕIUH,�	����	 ���
�C�%�k�9�Q5�w�.�����V�s��3ݑY�*-ߊ�'Aaw  H�e��	:�Џ֋*Su����L��_R�S!��0�_��z!z�Ŗn��DfŊ�㹵C����	�0���]�Թ�.�r��Κ��!��������[�6���s�KvQI6����z�O��n�i(��$��(����z(�jC�5�_�;R�b�y������Z���{����՗
e�Sw�ν�2�����UZ����_�2?ɤ�/��럺�S�}�/�3���[GL�|��7����֕�TDrX\�J��Ҁ����]����Y�@~�GzGD� ]�G��*u��E7aa�2\g�����V�H$
�/�<���B���`�?Fo
���Dxi��)c��4K�=9d~f�%ں� �;v���9	�<����Uj�(���y@�N����ގ��	
TJ?Z��/�H�so��@ܸc�Բ���	M�!��eW��E��h,$������nz�n�9r�:;���T��EOP,N6IGZ�+����;��c��Q�h`ߞ��Xݙ��rQ`i��*I��r�b��[7�7�G4t�7ǢR:hrͨ�����c�jd�Wa�3�vo���Ɲ��K�&~�$�'̩aBmN�(�<�2��l�����]�#�|7Q�{%`g0��C`1&�eT�i*&b©����Ӡ���:`7=iN��ۻ"=�_�`�U�3&����O�����95u���8�NY��%�kq�����+>3P.L���E���1{~�u���&�*�4K���D�ku1f��k=���
�y�XvD��
c��:���!��" g-ѡ�J��~̜�3���f�����A��z��w�#���L��,���:'I���xn�,���Bj����U
����Ӊ��T��2�L�۱���T�ʾ>���˱��4�vnw'���UK����}��wc�i�:��u\��-�3(�`'�us��>���t,�H1-�W��u�TF{oB���l�P��Α���6l+����^�.��vZB�IO|�((MG���BB�	�iȃ�\���ݏAPװ]�U-�S��#�tg����.�����i�O�!�[�>H������k�&6_�ᓀpf�.dP�aQ���}ڿ���9����kO@'�s�|�����-=�
�q���qt/'�"W����ǫUk�m�?&��z"P����N�����Y�~ϫ��������I�o��\���/��:�և��DOqyӟ�9�M�o����?������z>�Z9�?��}%RW�;&<`z�L�Ag��"V���O�,9	'h�3�� Y��s�F�e��><v�W5�z�} ��/����~��O�nI��Du+T���Y'��D�����%��9��T�OM�c��K�랦O���@Q�Ձsk��2�i׺}K��^������OW�� �ZG}qy_��_�eL�\��Mm �q��%��<j�3�'h	=P:����Cos,D9j嚶Ю0�r�6���dz�ŝ?6��T���#0�����O":�?��NS. 7/�r�Xx�'� �I��cT�VFH�HD�[��Y�� �`6�$�a�1G�+�����Ma%�
 ����i~�x��z�q�~t/���Dvѧ"މ_WE_f�EG\�VU�oeu��Q'����P4��:�^캵:R�h�2^q����n�)dԜU��M������7��\�7C &�EՉ��)yJ��{�૜��Pn��$Z��K齷V�_������zC.����Ma���mb=�}��������+��2���zr�sC��0�]��xq�h�:RSY�v�u�u3�]7�4$1��M-1}�:����s!3:2�Y)n�%o:88j����W%m4�d�6���INM��d�?!�{7�߲�Ȝw���E*�0XK��GmeZ������f,�}��S����D�G��]��K���C�3O�*�(C䮇ϲ�<�A�h���.����]���R�XB�e��g�^f/j�/��ㆄ��odޚ�������H���0�_���� i�3�/��e��sTDK��;V��D­�o�����Ab��U�����Fy�ԋ�i�&#�����m������%,��{�4/\8���7��"ʀ��Dh�	g�0t��}P(rJ�`,�+6��e���U�:��@ϡ�r7p�k�1o�n����� 	������n.��]E��Y�dT��D��±�vH��٣JҘ����j�@Y�|� 1ޜ�H�z�b�$�J�$�� =J���N�"K,ZQ�$0q�s��{�E���YH)���i�VI����o.�_26���B_�m[���jy�{fJD��&_�(L��4���\=�e�-����q�`9�F���HsT%I�//�G� �����ط�)B6Ϯ�}�񵄭�/\��+�����V��U�5�gd*������k%�>�����3_�r/u�(�HA�'R��-8��=��z+��Ο�B�;~{��Q<Q3Odl`��徃
}���g��l8�Aܬ�N��Կ[�`��!L�-�kv���v�1�|����\���c�������
h���=M ����� �ӯ� ���M`-B�^]�ˈT���J[�����3����d�nJ"��&�7��8����hvu�%c+E��+�~=ېŝ���I��
�|r[���Tw��$?���e�1�e��U�q7{蒄�vD���6;���rī�' ��W=*ζ�1�X!�Tw���e�YB}eg�|���2�j��d�%��S5�C?�P�gK�K6�7�x��|�>?<�S]��ƕ#�_0ђd��٪�!�_>ǎ��\?'W9~���c����;��ذ�ig��@Ná�Аr��/i�ZLl(����S���=�uȿ��1(F��i��UQ�]��H�7�b�qzt�4ݗ�^f���%'|@  ׏��y��l䷬��.��X���s�e~���]sښS (󺹪^X�#�� Ҍ����c�f���\ȯ�z����QQ�n����$G���Dz�59��>9s�]s��kv�L,��+̙FК�O���_�-� 
L[��]����9P��S*u�;,�D���g�3���v;�ɂ��D�������`�H}��B�Il�+�����7�j*����+��4�Yř��4�o~4`r>`���V �~���F��52�K���#>�sWUb��"����lٴ�|!�sF�.���[JB�'�u���nd�E'Q �\���J`x=���;ueܠ;mG��-�ry� *�I���v��<;��B�H�0;�!^)�2Fn���#/Fb�kfj��`��MطT'%`4 �%�kJ��ӝqZo��Z��0��rJ7�|SC�}!1��L?n���j����0g�N�z����  m�@Oh�	��q���HEw�����)����Ήa�ȓB��U�Q��Q��@���_i��)"�*�v�o[�M>.�׹aV+���!���W&Gb��Q7�	�Q֢����<�v��{m:�����ݕ���T��� ����78����b�;��-����a�X��74�>0����@c&Dh�6�9[�ʥH�D~�#1�G��E$��uӌ�ë�Eb��r�P�܂���Y簤�9�L��a����5�[7r��e+ٝt�	�&�͖I�_G'�J �q�!�u�D!]�%H���� ^n?ʟ�埨�D�#ߟt8�Գ�}0���T�inA�V���L��@GhFA�G;�b��d9~^\�]��KY�n�����jR�! 3Lr
ө��CXLX�$bb%}e�	Xuko|��]7�[�;Z�@J�)0�@�B#X
"B�\�!>��wv��,�+�
 +��{���[��>6�I"S8�D
C ;m�K�+u�J��נO��d����͢�I��.��P��^��?*뽞>`85#!��
�}��lEB##D_,�����|(�p��wQީd^g3Z�}�՗6f5=�پeq=�с�ST#$�~9%SF�e�j��6�V��I����hNQM��<���g��j�m�W� "fWi���M7�@/���F}����'�'�5��y���z���6'yl�#_֑h�1��Q�[ݫ��kp�a��K��4ٷ䰋u�
5k%�!"b�~n���)����`bb��P��������^j<�{^:c��*�V�B��A�p�����r�YZRؓ;pɃ��"6���G2 �W���2^�����zڊQ���l��<��X�d%h���H/�h�gUH��Y��>\� ��mCֽ� ��ҭ�-���p�W��d��p���O��N?��c���%~F# `b3Qg�����g�ʺ�<#�_��Xb�:�9��'�W�~�j�Q٨iJ��>̻)�Q₧kh1�: CXm��!�K��25�n��(+m���eGE��Llb���؅�ͱ/�nl�нx�6������I4��\	9������J^j9B ҙ���ތS��/�L�I,Ln�O��Nٻ}�JQ�I����7�H-��R����籓���Z�B�U�\�y^�z�t�������ˀ��!�M7��H���S$	��a��@G"d��=X'�+�]/(��\O���r�u�_N��c>�����΀��(l��9����4z>����xZ;����d]�fv$䢔��BQ��K�W	��`��g^r]Xz���PXN{]"���T��!2Z/��AJ���C8F�Vrn�KH�����ٖ��,Ռu��ŏ���M�Tf=�ԟ`jN��Bm���t����|����p�R=¶ni,*��Z��@#']��0���:O�Ά��Y5l�m��i3��Y	U^qp	����h�/��6�,Z����:CW~��BF��]0�.�?)�2���r�[��9�ԡH҈nLy�����V�d����ӌh+mE�JBY�2b8�^]����/w:��U��4v=�f.��Ѵ��	���k�lV�(��[�)�8��	���ڏ�<׽sX��-�2�C$�U�'VN#��s�o��<���*�����㏧��nݮ���޸|Fl����ܽ�wz�+ݞ.4���cv�z��^G/IGم�Z]ь�YPe���v�[��r?y����*�a21�����	��}�u�uQͻ�А?�+_Xs�ͯM�#/깩Y9W	t�n��/�;�XԊ�ZԖ�Р��Be�HBnv�=,e�
t����M�~v:�����`V�H��
�I�2��v?%dmu�D���O[��ɐs�
�5�d]�U��;ŕ�9���^J!4�K�k�Z�ix�n��#ũ��|�^ڐ)R�Y���K���L��>6�L��� (t<���@(�r]wA�~�&OgWB�&�/��FAN���0���O�����b�tlNx�e@�h&^�����I4 s2Y��S�4�,�h�`�����m�yU>����F�
��	^������s�I����:a��~m=D�	Gn�R��e����Ӗ3��=S=v@��:�zm�Mї�v+�������>�-��h�TU����}q�C�2���c._f�ҏ8lT�C4��bT^���⿼gi}�E����܄��̴��:[�	�H��s��-m�Y����fJff��UvQ��\^86��-����l���V��`�F��0�����`���ª9���>�N�1B8�_?T<\�^�d�س��z�MS�J�lJ�C�{
��ukK�d^)�+{�FϹ���*[��ŝr6IS:[����,̪ �Vy3j�]:����a�,��pp=
�����L�ſ��ϣg���35} �z9%z�@GN�s�޵Վ}u�聄����|\	�����P���Lβ�(.S��=�L�yX��a��1z��6�>� ��>����S�Oت�\3F-}rR��V�Ji��xrB����y���n�Aq�j�l~��|��b@6pQ�fc���vJo��\Hs:D��zI�Bq�@������\=p�멃���L@i�oma3"����	�����>���PtxԞ��΃��h�ө�n}P�D�\�t,�i��w��]mA�D��7>���)G�N�~y�n0���K�"�V�p`�p���k/��~za#�ޅ�~SI(���+HY�s���\V̗}
� �8w���zs��g�`��Ԝ�v���.�⛫&UE�>��8!��}��m������¨B�imr��S�*1$d�{e�s�c���r*-V�$��Y�ܧ�8��򪬏���7�	�o��E�H{,H����zF)�c�r�{��*�R�<�^Z������/� P�>���Gmj��˦��Fքm���;�{a��
l���5�BY��I�h��4~xr��	��w�$C3 .�ອ�-L�ظ[.m��=80�"j@���[P�� �K�X�&m�v
��мV�<��M�����(�T��c`�l% n �_z%��G��������e'�I�V���qC��s��l`�df���7��n[����I��#���B>�s$�_�s��3�	�O��{2�(L�hgث7��$@JC��9~��QC�/gb��υb��:\��q���U��}GhQsW�B�sZLd�LhB% ��"~�7x[��Q�
*�\��Z��q���ؕ~Ӡ(�.~���ڮ�zC����1���t㨔�8_��r'��[1���{�c)�f?����g4�ۻp�n���-m׀��4��[�iCO�L�����a|��%��b��������On��;ӣ�7�p�Ϸ�c�D���
b{�	���2me+�@�ɒ�o�yG��}��j�b�4�vx���ƍ|��łi��%���N8E���]�ɭ��[:*VH��#��z�����=��lrIxٔ\��R���T|�ʲ��{��?Q0��D����3�g����!^:'�N��:����-O��� ���5ӱ�%nȧ���y�-+���+�"�qˎ%�o��ޏ9J��Ig��D���r�!�J6�p7�㺥����37��ĩ���������^.��,hC��Vy���pk6�D� �7V��N���U��`��3b�$�,�w]o���Ww8�v�\?�B!ٝ��<���r^֧�і�E�^^
ۂ�=�!�~���[΅1��G���Pw�p���Q�+;M�ML�"�:t#}��ـ��*��ǎÿE��89���'�L�ï�}�|7C������0QgT���)�ʪ���-�~�p�z�?��J����t.h߸��V��J�j�=���>�e��ב)�WZ[��ʼ1"g����y5������ZZ@aa��;zUo��/��S�3�0�������.��Rw��u�q���R�c@N��i�?��9!�)-�H�J�Wt(������gE��Q֣�+l\+��txP�i2��!���'���q��/g3�����T���zl����z�ab�f�����%���xT��|��6�;���JGs���$�#W��L��/R��/e��4���
�����?b����� P��Q#��Zc,DxQ������Yv���;�R�{�u�} ���՘ͻ�᪅��Ċ�}F�� U[O��*@D~+�П�����[�SQ��ʋCsE]�Q���@��Ǯ��/��x2���Y��e���X�L*n��}B@
�:����l8�m0���B�-F�:_�D�E�t<kBN���tRN���S
H��CBI�ľ�����v�����u=�l�3�iص
q+�1f���z�h�"�Ql�,���g���h�vh����_fqi� A���2'�t�w��
���I׷��܆��F�P��Qte5����;��nUT���cs���ڼg����t���T}o_rە�Do�&�'�r�������vK��d��FNDʕ��ˇ�%JJ����=�w.�;��X!�?1�9�v8S�b�57̐Y���/s��*�ސ�J �<�[���`Z������T�����+�3�[��֕�_�a�-��!��Z�;H��p�^��y�V�]N���w߭�}�ķ��]v1Y�M>�et���n��e�-⥿mG�y{�@	��拾'@*^�F������\۟�Y�|�G��{�C��BK��M��WM`~?w�ki3헙e�׷:W�z���B��sD��Z�!�	��mj���V�|�J�k�c*���
l8���B��9�cTV�öRt�����9G�����*�f��l�0⫁�e:�[<|QWG�6����@�)��jҵ�7�"Mp�Ut�n�e�+H�""җs>2���~����%2�_�=��tV�/@&u��9��ҹ�8����6�VX4�ڶ�&m"��P�����-�~����uB	�Zr�p��s	�%��_�#�?���|�8'��U���b����2��UF�7kk�/�D27_n������z�=̰H��������w[��B�������S����.J�M;�p<���rtj�v��2�I��I��+�;Ӷ�5�/ِ�Ľ�g�TF�����v$��>}n`rYv=�(�y���-[��u�w���i������NU��G�@�G��~��1�NyQ`}��dAu�,�D��d޷ E�J�*V�I���$�ń����hSmVT��N�Ƣ���M�U֨��������Y'�R���A�@��K���7� 	>f���B���69�(�aK����-�I����)ϫ����bX<���宥Z�����������E�^��K����Z�%�1�<h�ښ����42q5�B�i�D�ܤfm�sw �����oo���*�@��\�)� �/H�����pI���̇�6�(EHOW
�m�N�=4�ND،�fW� ��4�%�с��)�Q�Ý%�N�����*[��t��y�6?�/�!�r���tPX��*�*�S��ޕv��Xe���>�e����m�?[�\��s��8L�SZ��^��V��T��aJ!�C\���
lm�;��=Aa��W ~g�	�9B$���%6��!zغY�U�n c1Sȝ��̺��>���I�V�2�+�&�"��?����)3��)l}���Z��χ���͊X�D����I1Z*��;�5���\@�T��,X�e�UE
�izxȋ!x�0aLa��t/��>�Xz�e�)�-E�_tx�~���4�%Wc�]Rp@g� ���(�Eb�o��`��:?�[
 [	�e@oʺ�h��Dۿa�m�N`�������?�~qm�5��Y�D�_���E��;3�4���N�ڹ��x:�ʚ����|º� %����������7m�e� ���5"�n-_�(yK��W�W��9G�
U�R�|6����T�ls�����"�(3���-��h��vIN�d�XtX"�K
b
LDH���K5��pn{.����Ão%�OV��)�[w[���yAv&q3�'٬�w{t�̞5���� ���[����Ȫ>�y"�׻h��t�'��.0IW ���D1NE�,�(1ʼ�����-sF)����p����FzD]�LV���|>�4�jI�f�U��)���͙n53�b#���'�B�?�T��lzi���5�턊:�~��y�N>l)����?�1q_! A��I�@��5F*��.]����g�*�E��	�S� �M��NS�ܛ��T�7;�A���gs��G��+����r1��)ꌵo	+��ba����;�N�CA�=�Nu.�oo�լ�Ϝn�$�r&��r!o͝���Ȏrҡ&y�]T(�/d���cb�8�w[����"��	��G��_�����8$D��zD�ͼ>%F����r��I��d�u�gҘ�[��߭ ���O�y�k<�2��냟ĵ���yIUk�t����z�̫�|$��L$$}/�<h]� ��Џ>q'�~f���2[��o��S8��Vڂz�w!MIrl�]�D�o{�=�\O�ʊ+"h�t�V���8�ҎXGs~C�BQ�E����{����:CJ�:Zv����VдP���L����ջ���񉈸��2�s��>9�`���W4�m1���C!��3 ��8u��b�o�h>ͤ�#��*�6�A�Rc;��Hz�����0���^�ۅ3�.|�}��U��@��k�z��~�Ŵ��פ���{�Om��Q1"!Z�U��l��y���*j;�	s����f?ᷧ�g�����0Zok1D��r.I�����ܱ<T����&���\_��
7�tj�����H�ڛY�����M�!�obzZD\�DI����g9���?� mV2GX�աx�vmӸ��$B��^t1+��EIk>|T�S�}P�/�J�\݉�e��]O�	��g��9[��Z�d}%�����
�w�%F�f#��fC.�������_Ѳk�Ul���4��~��C�9�|�e�fb�UN�iT6�^��q�×܅� ��Np	���m�WI���;䃦K�^N��7�)�F�o��Bi��"��/{� '<(���N���1Ԕ�8q�?�5q�Io &|���T�� Fx��B��pME�{M���n":����c��%��_�T�����-�d�
G�� �Z�g��f`��"�r5�����V)��m�n����.to7iI���bH��l��M~�����AE�P�"�*�M�ҁ�|��"B�~�T$cC������d�����4[�7���҉��X��~XCj��a�h��ᭃA���xv��ӎ.o��+��ew��|��;�4��*˛�������y^)XlN�Y�^dm9��y{e�������}���@���&Wߏ�qŹ��l��A��T\�I���Ø��ـ����xZ_'��ʢa����|�T6��W&J�H����\���eX�1@��`x�_�*�t�2�21t��Q��h���ô���o�v���C�'΅_j:�5δ ������es������j@�Q�vd�y�u ��t�q.���o�A�h}ҴV&��h�3� ���""����5�0E�(N?�	@�H�|�>a1��M�J1���왥r9�s��j����Yc���Wˋ�3�.x��}�}��Y���j�ɝ��5J��$��%N$����8�;���S���b��
��"۲#u�9��cSV�ٴ��5��`^�Δ�|Q��ōǥ3i���
�3_�,��E�D� �1Q����x�T�{�sq�}$"D �x*����������c�ťZ�݇e����Y�w��_A2GG��]@�R�cn��~8ҵ�!e���M�e+�;܏�&�F5Ez����gDU���4ƅ�P؎�8 �[�gW�6h�c"k���(�����{�-�.�T�ŋ7	_�7	���v9���y@�|���^I���Ck��oZ\�q�D�o1n!d���W�^S鑢T�j�)�i��G�w��\*}�(b ^�|�×��n���=��k�2�
���M^-b�^�3"���"����`�G��<�J6�{К�HX;B\���[k�&���K�{�b�R��'v��-_FK�ѽB&����ۜ���c'Z��jԊ����jԊ��R TrUO�P��H�� �-�������oz/�,���c����T�p⯥\�vB̬4��'K�}Y5�����{Ave��;�i�Z"^�O����}�������Q���jnǽ
d?��To����z��򁟡���
\�-�����(�ַ���@��T|=751��[Z����,��A���Ȫ��ף|P��CŢ�o�\���^�Al�`�'#�[��ݲ��{y$���'�
ŵ�D��Y��E�O�'lW��+c�Ǔ��o�;)�R�Ë�z�5CC�M�Ê��8-ҵq��Y`��d�b}�N��)`��j&�b0�?#��	y�բ���8o7f�ߚ��̦��$��i�����L�3��*'u��o:�d��2�Sv����u,x\Y�l�h��ڸ�z����Yi�����(�6��]���W+p���)t���x�s��ܛn�n��w����Y�g��Xe)�fJ�z�=J�=\��D��/0_��T������㝯��@A�6k��^n��ۨz������I�l� ���ߛ����� ��B��䷶g����0���NoT�P�B<���:�1~VЭ��ԼÐ4n�!u#��S"V��:�k3^��Ǣ��Ƣ����]��ޡK��R�p������h�-��nG�����]�#J'���*�X��,���~=
����q����Z��xk����y��O"{�z�8g=m5l�Y�R�0�B{�ڂJ���3ni{��k���������z]�o�(���-�ԥ��r���&�nʫ�{��]�fJ���R�0�~�^�������)��M$����&�R�
�8lhs��)�l���+R0/�Y��������7cӑ��z�/���mIY��������&#����>R�O���

�Es��	ͤ��Q���r~ژ����X��S�M�lF}�� 1��]�n���!�� ��1/|�r^���[��� ú�6_h��T���v*�C'?�_����9T쟹���؟\O�����
� �J��
j=V�q�JU?�V-7.Q�BJ{7ud.��m(��l���Z��O/z���6��5�jc���I!�"AL��]�s�s���Jk�"�w��	7H?��ysqY�5Gh�;�[��H�[�6P�2kq�H��{�u:��_�1�آ�:�u��y�3��1�h>k�?U4} �A�h,A���l�3�?�A����'{�'���n�̏�z�ʗ;��F?�z8�`-�ש����u)Q����!f)?r���G2�)���b�$bڀE�K���vl3H؞�$E�y���Ǘ�EF�2�;�^S�/�Wjض,�i�!��N�rVMʺ��+��<��� ����mRHyѠ��YY��p�u��a~�,�њ6�U�>��9��ݼ���-}��h�O��k��M��?�ve�ܼ�! `e�\�:�)W�~�8��I���zǂg�KKVᩦ;����賲2��[�V��ط��	[jLM3����0�a%٢ϭ�JT���X�{��%�����
��ϯBh�n�rAj�S�==!�<����!�Vġ�b�#�;��<���6���R�3���"���F��f��н��wc��jGdXiT\[J��7�?��90����ɑfptS��U�$����\n�s��<(IH	�F8C�O<]QQ`ePG-���t�����?�n�9�e��s�F&���a�'����/l�:~}��bm�	�~�����^�muc��L�� z��#����|5�vy�"�X���w�V���< ���jD��	u �W#���龁j��3��)>?�W��լ,{���^XKx�<�*�^�zC�	x�n��ʮ�4*|�j��]�y�h�*��41Ū��`����ث�#�vȺg��d�)����~W�3��i�B���^<mZQyҬRѿ�2
���b���Ք����a�}ބE�����K�V;��bi� #�=�HX�-94���3L��o/>^C��j��_��Sc��Pͽח��5W���kio*��F��ҕ<����A���E���R�	�í:�tZN?�-���QNh�0ߺzc�t�a��a�'{�V�D ���Ƨ~�?�_��}v:ͳ/��x�l����9 � H���g�%��]_{t�B\�}�jKL~	��-���S���DAi7�=J�q��4�L��1n�+N("�b!���AN��u�e]Y_K����R#&�hx3\) �,�Q �[qT~��_�/��	�{�s�������-r�dn�5@��I�b4��������L�E����R�g�~�Vo���� {tP5���%$�����^�+����{0ݫ�G߬�i����$	�~7��
�E��Iy��d�07������Lw��A_e�}���/kub�������1���̝呀-=v1^`������������X|51���j��}z�U�7P���1ߧ�!��*����P��첤�Iv ?�� GH�;,�,	
R!�0�~\�ꎠz� )��n�;�_W|
����N[f.��M�;���%sN���;�9ժ"6�ǿ�N�f�i[Ym��v�,�=Bwb�'|(ܟ���tU�(�t�|L�������-��+����⡺�{\��$�3a��}����1�V����g��r^�������f��^t��"�c��#���3�h6I+)���ɑ���	J��f��O�+r��c�8z�t��B�kdY_R�6#�}����8�P��fN����X�S+���[�݃ʯo7ˮa˽Dl��0�g�ʘ9�;v2~�#]]�o���q��ܲ�n��SJ� �u1P�Ts����w,4y��G�|��q�E�(�	��A�,�������M��
;�̤,J�ԁ�'��dHO�x��U���/vޚ���:H0�����G�M�a�l���� �)�8	j�s��-I�-�.%��ߓ �8�1�&���O91�m	*S��s4L���j�I�s}IAv��^鴷b%�_@A��Ϣx���2����W����z4�d�j���T��+����O�@/�M�⣚�����B{��D|�"��S��d���a|� �;d�k@�ߪRux%w�ޣ$���5_��<��-8�����_^�kzt��i+���>�]$߸�sv���Q���d���{�汳h���LF�?J� �������
}ҙ[��b���"&�:7g�O �fp�Б���]��c_��5��q$`�0/!�A��=�S ��% KO�^�VE9~(�#��	oҏ8�˞�sI�C;��v5�y���x�I6��y�*P�{��Cn�@X��J������쏠>��g*�س�/~��a@�ó���*�'��L���b�g>�>y�j�>�^x[��z�Y�,��թ��[�6����Ԍ��m y>���4O�ǕZ���� U�������Y����F�1���6�Q��͆�)�ɗ��~H��'��f=Ǆ�ӿ_x�����p�$�z�eL��2fן��ٸ�J/@X�
Bx?$��N��g���!�}���i�M)t8U�(��^��Ͼ�㯴��|
vT^r��!�������۝/����>�������������IK��Tq6C������C�^���?h��=��3uchQ�rS�~�U��~��K�3�ۮ�L��X)���VIZ�"���C��☿�x��@��-�� ��7?Ջ��Z�\��}1��U�9�I��V�d��n��4��HD�	Ћ�p�Kzs}��i���aXd?��\D�j/�U�;�5q�mSg�����_Pi!TB{���_�@��{#F��V^��� �c0P_vc��^ea�lWȣ��W�;�z�Jb��7j�� ��_�f�ׯ�#�n�	�8�ǐ����p�]٣�j�(��Eٝ�|�4��8Kr�����S��eJ@�&p呿BթMVK���m�������~H�oU�ھcz�~�	�'3Ё�f��!
�d�sb�X����
픈)�L�aw	�DMϰ�a�A�<8�2�k��"�ws�F�du�����;����E%���O�i���_(�=Ԝ.>��|�c+Y ��E��R�k}a ���PB>�|��
���bR��P�z�)?9g;1���r�H����
��܂������ݙ����A·a�n���ֺ0�Ĕ!�GL��(KcςA�S�ȩňR\�yY�_��G��8#��9��i�ӕ�����G���	�ƪ���t��sm��A@���S�+.�	R�FƻDך]��z �E��2�8ҩ��Z��B�_Х��H����@�Γ*D���&r)R�{����T�_�cV�Y��T��q-(��� ��DzP�I��t)���k���B�t,)�jP:������~>���7w�̜�+sgg���ma�i �Tk�ɮ�����аu��9`lo��/�9n�{�\%ċ̩�L��;W�6h�P{��&��,+�PN�!���ɽ2��͝�����S���Ņ_o6�W>�^��ڮ�Rқmp"����_���걺(s{����%μ�=Ӆ�k�'�oP�����Uh<�m��mi��D���6b�J��Ȇ��,\�	����	��X%���W�l1�y3n�a6\u/t
���nx_j>-�2E�����=�*FuM{�lS��j�0z�|x�	�(���Ő�nGe%eph��}]v��w����&�}���oK�X� ��:��܁e��(����ZAT���
+��� }9צAT���;�An��G�x����7|u��
�g�E���]!��9�}u�	M����ɬo���~����'��E�����z��#�n������6G��^ͳ�� 䋇�0�q`x�w�b�!���dV�����CŨ�kk��Z�*2���G=�ש�]����;LVd:J>z���x!ס�%q���3���)/R<�"���(]JI��f��o�Ny�1��~�ވ���B������������v�~h.���AT��Fr ���2Vx�Щ!bIK��<�Z~�刧@����C>t'C.P1�9��tsfY^�ѥQw_������'��Q��zD��~���~#�I��/}�kO�d���j�=d`�(�bn�ˎ��!��~���9t��M�)o�0@'���l�sq�j1��@D7ᒥ��Ѻ����5� ��niOirӹt�*���fcrz�gr�5x;bU������;t�z��ջ�e^�Xf �#sH�|w�qxL��0�O|6 8U����C��8K <�7�8��p�d�$�d�<0��{+6F�:PZ��b��s*;�A���"uș�h`��(vV��'����e���$q �	�?iY���l���F�>����ymΡtb7s���j՛5�Rʡ!J�y (��@ݣ�p"Bi���A��J��g������-��MW���'�\�� �N�M�vm]qBa?���EZ����$0�JHPF#s�Y�<)4��ǁ&�ӓ�Q��e�ա��˶%b�Ċ|?��h)���7sC��㕂�X"��g��w)���t��i

�i���)r�1��x*&����X�I��<Jw��Z	�U�;R������>Q�=Ӂ�h�¬��*j���c�y�+}�}0'��\�H��e�t�ic!�¬��R3��p]I :i���zms��z�&�K�g���j�z�J���Z͝��UW���19<$�ɯ���a��,�hiqgj���
��(��s��Q�&b;R�N4p�,������_}8\:=�yI�ۜ�P m>�\�9��&(���]���7c(i�MAF>��t��?L�x�ut$�ji�1��鼔ה���%AN[sP��a2��?11�	R4I���-N%��ڥ]���*�˿�Ū����pһ�t�D��Ǘ�!ǉ�㴔����*y�����l�i��{���D<� :g�4�MM������5�oo���ݨ�΄��d�b��F�����|�+u6��fq��w��'�a�����6%��!$m��(���	K�X^٨�	 �������c�n-�����y�IfsOk�GI�g�ʮ�O"�9�4�����\� �H��f�N���H(h�	g6�ʹh�/��c�mG�U���a�⑛�mYG&/E7OOfQQ��]�:B����'S��'�]�o3	��Р�������6���d���g��D���~#o�ת�J�L�΄��6��A��4�$س,!-Jb_N��jl�@3�5�A^�S1\Z��Bx���>�u�"�z��G]�9�����[�8��hC��f�01�U�֦1 �3�C W�̉�N.Q��kR�^�&�o��1�6�#X		�4�-�v)p��ϭ"^���d�.�Tc��W8"�h�ۏ�6�2�۬{�%xmH��H��GGz/'��4�c�*4�T7.'e.ѿRmivM�1�k8��{q�n;?���9/z.�l�Ɠ��m'�]�[�EHA�եo� f��(�jN���V ���o���(`z�{߮/���4訕��>C�;�i2�i��K�Cݸ�s�������Sn���{]�ƍ匛��=M��R��bs�����cz��U�%t��Q�r�܊I���o�z���'��.���VJ wvԽ���=���J&�ӎ�܄�(���0�@�1XͅA�К���Q�R�&A��Άu��G;�K�2i����)S������7e��%)7��6�<���i�Pzy���,e�'cz�Ub�!�k>+�3M�1��j;Q���Zsw�=*<�y�R�o�jv~{4�4JWO5��Fr䬤�ZV���y+�"����fB1y��G�W�eגk	j�%Eh�}�Z8W�u�]��XB#rq���J���1r[?�:��6�m)|X���s�/�O�����M-���7��Ӻ��n?���pIW��3ߚd�o;��	�d$x��w�*�Rj�_J�~-�ZY��*�vݛ��j�k.��ʲ:��L�YΉ˥@^ƴM���S˝�Cm��B���0�����M`fPU�@D��I�d������i��2��Qĭ#3x��CD>"
�����p���gr�s-���EI���z��}[��s��4l�<�5���#�u��Zl����<�q)��`���GV�C5���N(���|7��S8�I���Ƀڛ`�Ԯ��T�]��I? ʇ�i��r�5e�넺��J��LT�����B� 7�S���=��.�]���ϕ(gc����.�e;�D�*�m0~x]��5�>.�nk��aa�?%>!�ډ�������]Q��'_w3��k��C^6�Y\ Uf��y���ϑ~�d�6��z���*#��M�u9E�^��[��ѷm�0Hc��n]P	�⭪�4��h_�dcb��{�НնFGU��a�}0��:����Fs}1~`��-��/�S�|��� ���� ��=3塺;jȣ��mpH��і{v�\���;�Y\���c��߃e'!w�w-k�5�nѰϏ<�
 O�{A]p���j3ָ�hZ��^�u�V�eI�f�̛��R}E���Bk�Û*�,���\�/PD����F���#}`j�����	Z�"�G�an3��
�'�r`������sU.[�t�!!(9c�铯]�����fb"��l<�~֏�4#����೵2~�mg�ok�K����/��ds���gq�^�M��窊�.`���{��	�k��O�绑�D'v��ߗ3����7j"J��0�K}\{/:Ӌ���ۄ��n;�����|��zx�C�T����.�A&���KO7(���_�wJ�=I}Z3*T��h�����,�ssb����R?��cG��?%U�L� ,,
�"{zT�(����.��`b���|l�A7��q}(��4��ͻA}�ќ|%nXra.B�v�ikC�,�lӊ�j��ى�\���kԵf��}��]�J+��k~A�+�U5eG��Y��mPam1i�<=��­����G)+0������+:A����R��m��3E>��zP*�����U<��w�5�~dg �nz�:BF�S�ݿ����,]=�?���Gv<a�oC)��%9���ujC#D��8�dʹ	� ��{ ƥ=���a$i\{���^;�x%�0n{����G���Z����K�4`7P��{?�,�� /��z�5�b4)۹)��{U��f�A���{>��G;��f�3l��B���E n?FT�Y��Y�p��*�6�6*T *�tmw�X=���x��ʋ~g���C3G�����.�q�lK�X�շ���xKo=6ْ�Y��2_���Φ�E��d��k,|xb���+��H�튚��N)��{t%Iq��_9�J&��Q�������{1�R�����D�@ݲ��6�7s�Ŗ�o�����-���)����7�Y��%_��B��x!W��F^..4���ř�z#�*�r��b��äT{�͜i��˩���I=��^I��R����+�����&t��[���wv6ˏ�8	#u����L(n��o���x��^�}O�E,���W]�~�@,���>��TPr�3�a�Cf�CtRThg�t����1���LĢw�O?`��ۣvY�� (-/�h��;&��P�ٮ}��� gW׬/?�-��۞F·���6�~�������[.�ud��'�؈p�4,��W,0rm|Mo��R�8��_���9�
�|�N���SM� N)T-o!i!U�Wv�*��]`�c�l4�ic��+y&�S�J��6�TD��7�^��OMSj����O�S� *�H2dcW�7��DHy����eI�G�1?�����t������?��)��1}U��e���{pL⛝W+�z�Z���5������t/@v�[�[�=FK�[3�%Ue�:vg^D��F�#G�ILl�k��E,W�/\ka'}+���_�{�)�L��<��KW��m~�!p��kʓ��5��Fj��}g(��.����P%���n$��̊�O5���ോ�?�z��	��O5K������L}zF�ݯm/�H��G��l�:ǥ���- �y7�u{�l��ko����p�Y�?9�o�s�W��n\�TYqQ:�y��A�y���!�,j5�ٵX�'h7����������]X�
�^Dqֱ�^�VLVH��H/c�sn�5��'�1Tޠ�lw��H��TI���b�̲*��R����._�)��AJ轥Zˈ�ZЙ��:���K7\V}5嘖���+}=Vq%�Xh}:�b{����w�'bb�_�mo��+d`Ž���6%o�F�m�V)[�fkO@:��<�&�3;��֒��c;�M��DzB�a�07:�`�N�.�Ҽ�����.ٝ�+�"#��d�ەںe�����R8ѱ,ꦓr^x폫�xz�"[O��Ӈ�y��&X��' �)�"q]+E��SM�q!k��f����)�]�Jc��¿�v���K����6�̾���(.��;.��ly/p{/�w�d���y'R�-l�b��|C/{:���u���^a���}�?p���J1����F��˧�v��:P5z���"wى�%�F�	�� �YА��ʽb����q����W���+�X?�|t�� �ڂ%F�H.FF���[��]�BU��/�M��������o��������hM�n�&l4�Aj'��HY���;���2{V��V�7o��(z�je�5�1�M)i0X ۸�I	�W�#�R�_r"�����F뮷Q���3�U�7��j�-/	��Ayej?�������d��I��P@@�W�'42�0y#��J�{Fq����w�[oa}�
Hk��>4F�+.�b�v�	*�v�f>)��b��*�sSUt�z�ʪ�*��b� @����	f�ZSp�^֧��]Yq�����N
y�F%>�[�� ΢��kØ�Q��b��IEv��Q;/�d�!/b<+�zk�	�
�[�ڑȠ�Qi~h���o��=f�D�Ӟa,�Bx?���e�7��v9ᙴ]Fd�<(��o��8�}�EA�|��ݫ��>抦��N�c�6��AM�v�q�cT�J�=�rU��z�v��^BQ��h�Ni�{lf���?~~e�`#�Ԧv;�WIv� �=�BΕK&�t�<Su����4<�Z���䡅JfC���O����}{��/����u�5�E��0�}Y���wjV��,.�|n4���g�,�e�=��)Ƒ��d���ȃY84k��0��#�A���.��Tg٣�(����s`_����$�\ ʾ��j�>^�/���+y����es輿�zЯ3,+�J;����QVw�@�:�C����nB��X�W���|d&*��9����mE	�p"?�P7.f]3Q�t
ۙ��-�vb�&W�;�����ixL���[�1~s"e{�����{�Ew��w3��
vt|6�˨SL*���>A��З�� �l Ԧ>�q��7"_��.�,�O#<,M�N�?ag�Fj�]�Q���ݣ��c�3Rޔ���>��I��饼WW��� ؅%���Z�t����/��(�4�Ķ{�c����S=}z#�Ǩ�"�A�`��8��tޚ������\N=p����]z:�Z9����x�Wc�V>LeNc������P+7����T��ڱ9�`�s�f1����H�jlQIV� ����>�g����Eg�j�CAX���\J�,�#�1�vЗ�,�ߵ]�,�<4���ݜ`?��gLl�"9�}t�A�e-Mu|h�UL�'�ϰIR�����K����i��b?Ǧ� 7�U��=�HP�������"2ϗ.;ӟb��� =�R�r	��<]��c(J�n6��Z�=��X�U�[���9|�7Z��x����ɾ����*��}���r/c��ն3�<$o�IO�Ib''�<�O�˽6�H}�H��$���%]�=0�T�9��� #���_����m��	��o���K��E�]�`p �0���a��Ny��#vQ�����Q���#�}ɛ�f�0g�赫����R��s�&<�]�k��'6t=`T��WJ+��9��I���_F��^�����|AuJ-�W��Z�ع����fB��JX?�����]x�A���Q�~.�e��5[Y5��QQ5�����y��õ �d\B>RX�"X��,��/����9�O�Ur�*�$_�)���x��֫���j�#���yu�rT�t���w�3��BmhҊΩh�%B4G��8q:�8e|U:�K1�oN?�X4G	V.XbV,�o��;�č�q�ot���W㪈u��#�JT�z��ި��8"�{G���j�Y�?�~�Vw�S��*�mOKUy6u��F�<(-}���j���0�R���Pc;��ٌ�}pήg8��K��r�'�Б��D���h9�ta��)-*-s:'*�5~U9F6���d՗�P1Puxs����o�/�H(f�������ր������< ��e��<���sA�PxR���=)��Y	�f#X�U����6����BK�[bA��+���M�.���}d=����hNd~8�軆v�|��V����e�J&�4���". x>�1�
H�"�P��!������]˗��t���w���;��Q�Xw\����7]�[o�ɤ���B���4��MN�Sw�΅��i�u���彧Z�E&���U��	L����n��G;-�f�WQN����; Nj�E�P?���{��?�ON?D�-b/�<K��ɟ֡��8R�gC�����a��y�׋��8!����vo���z��,�
�R�}P酻k��s����~F��]�۪H(���n� E��>�S!�8�h^ *(��v?	r��&�M�K���H ���V6�b	
ք|��������N9���d*�wCg^�v"�6G�kN�0�5�F|��&6y�w[����&V7;�c�:r�*e[���h���F�_��mM��=��cW��$�����W��R�~Ȱ�3?h�������k���I��<M���Q!!�2�k)R�i��������Vp�j��=��WRL	�zX�لT ]�m�Z��LyM��J��Z�Eɂ�~~(R�o��)(0n�v�9��77yU�G�>3�]� �Zj�ػu�U�8�����iP���G;G��r����&�MefM�N<e��SM�u��]>t�����;6y��bDo\ �R���bc%�b��+���>|�k�76(7�����]��W���hs*��.�q0008z��I_����e9�,��-��9i�37��m.� �@�'���0�m�MS�er�ԕ+/a�������N_����/��
l�kœQ3I�^���Rv��d?t���x*�oi���w�ҝ;U�;����5�.����^O�u9+�%|���T�fd)��7�7�[�i�J���$`���y����x�Mwж�hX0�Q�Jp��x��4��Ɛv=��d��6��ݍN��c�~3Q�dz0';m��l�W!��aO��\��*��a�ȗ��$�_p~�,�Ǫ�q�*�����p�ϕ�Z���'����*���ZuoN�iܾ7h�gr��=�^9դ�ʼ`3>Y�"�R������{���c-��qoDġ��L�n~ؔx��@��j�d�����zm;�j2�݌vd��Z�"���9����ߨw�ef��ȼr+h�W�b��+�n���MH�F��\h[�O��;
_�`�(6����~�n�t�B�P�4�<˚s@~�cC�;"���cX@�ռ�'�P�C��clh���Fg���5��ψ�f(���/�9��G�q}��K/�C�kR����=�͞:ޒB�%�-�aƔ�tM% 4��D�_7�x^*�Y��K�ڧU�q��?�`03�o�8?z��Im�w�Df�ƭ!��QA��浶>7��1�i��5#+vl��Sor
?(��<(����S�z�2��5�#��B^���,���V,�~�N�~�u�,y��;��TV��Z۪��P�;�u��f��޽���1�h�F@a1{�l��[d�-g��? U��;���n=w�rk:V;�����7>�uS"0,ƨ�a;O'>guz����Z���O�j6|\�m�\�:����oAv�������+ZH����3��-T%��8�׵Tލ1�n���Mx<�0��j��/N`u�z�*_V�ap*	���)���4��;��`<{��+��o�R��g�}�7�6(K��ě��;;�+	Ǉ5�tKC�E�7J�#!�Ү�b�i��Vʱ�|�Œ�RE��QOL�K`��ڷ���$:� �}�\thR���S�c�n��)#�?�芵��h5]�g�\sv�!KsX_��Q�L�K��'�u�z
.ٶ�zA��D�|�����#ѡ$t��k�I����8DF-!h+��|�B	kk�G����|^é��]o�[���V=�|���\J3� u�}sn������@!;��lш�z��7?$�3�A�_�rC��qB,+c��}7j�Y�{���|ӳ%�U݌��#�>��K|���B�H{��變��E;�[�h���Y��:H @呓�gt�=$�\��c�DOx�P�����R"���t�o��|U�EWn�t�%ߟM��<#yfiV����[����^[���ZKY~n��<�t���^<�3�Zݹ��n7�θ�MU�|�G̹(�{{4mk^�ڮ����9CT�`lmeO�����=s��0`n�<�ߥz�.~�E�O��뵔?�c��q{�)��$�y_��ȅQ�5�8얘��]� <"���>?I{6�(k}�hPS�̣/�$�����jrZK�d��-'��1�š��`�9U�U��;�+�'�ۆ�X��Ee�<a�ɏ!�*4ZT�9i}J�d��G#�.��-s�a���h\wIP�O[�(�O��**�Ox�]Pʾ�RZ���{��k�dO��>��6s�^^�Y[�;�ކ6�"�I��33\�k�(�jϬ�׵��%��)�ԯɩ��9"���_�e2:&�N�K�>���P{k`J��	��e��[�U#�{�<S��������c���L�'�1�`��߅TeVVֈv������O}3�9��i��ݦ�zźN��]�\zQ�[�ԑ
����2�p��K�����m��>��#����Ǽ��p�y��i�P��̜�y���9������[�7�S%�o��|��nl�O�=1�rX��jﬥs�dN���B�
�@p��v���\��1��se�$��-,<� 1N�qs�{߈x��/��Qa$irDkߩ�m�o���y�ɰR�M�Gilě�b�k��D�Q����;N�.�n�uQ���I�\��=�3��be�����3݉UǶF�����59Sϯ�;3�Z�y�����}�q�o)����<HH��w(Z��O6������q�cf��}O6
MVHd-e ��5r������\�p�y��yGt=J=�k�v�.B��!>d�<Ē��|�#�`ͶLĆ�u�[o�V0�s�����=�A�F]��̹T������],�C�����=��P���N5�:�y�g�[G�QR%&6l�Mݫ)�Yr�z_A0�Yw/xՈ�Y;��e���f���4�<�e���p<�'9eW��E�m���\���͝�HI�1�)Q�!>��g�]09���|���kw}-^�-���vZ�Se���� )����B��ٯ�F�^E7ښ!D�W/bi�����q3���$���b����.���Qʆ�w�5�}hZ��VͿ���pmx�����;��J�����6=��n6��m �Г�d��o����I\0��%�[ڦb :s���+������|J�hj���%h�Y�O��:�����ߊx����=�Z��+�x��O�o����g��5��u���渲`5'�%����I�)���Kځ�-
��LGo��	^�Si�~a�3�^AzZD���Þ�"�&��wN��[�>�E�'x���]�Y=��"�!۬�J�_�L��15X�;�[y�B~���P�~�D��;wT�S�*���H��1��T�1\*S����t�L�vvmj���+(OD[�o9��U�z��i]Y�2��9h�V`mN�奒��k��ȧ�{*}P��4jh�`�����Z���D�pQ�s"�ć��.�n:�n&a��V���435�<�(������i9�� /��yD�l�j
"-�CfZ�o^�ߜر�j���p����o|c����{�.Ъ����։�y�&���1���r���7Cf��g��Ĝ��dK���̴]AU�6��kvW�?�'���фv- $wB%�.��J�����!u�7�~�� �Oi��L,�9'@"�˝�H7�����/]N}�6a��?�*�j���i~fiQ�Ҭ��kD�8/����&̹�Zp�� P�y�|�8q�p�̒i��o~����.��1�q�$�T�_����>�òk��l�v�R�W>�ab�CT���Z/i�� EH�h�Y��*DQXH�0O�$��=����.��;��/M��kW�׍l$��S�\H�`��I�, �0Î�+��.s���1�v�b��{�]|�ͺ_�x�-��GE��d��+��*e���U�Mk���������9�+�&F9ʮ(Ä���yy�<���?x�q�E�^o�n=��}�Dۺ���n"-)�'���\4(5���%��,l�˰�~�ڷn�p���u��^�p�Wો.�@6�����9��Q��ӊ�PfZ�i)WL�2Ϲ﵏k�{�����-Z����`�L�*FGB��uz���uu��nhe-�S�;H�\O���N�]k��r�o`8J�,O�����K��
z���h�,������4+�x"���W���Y�>O˹*|��G��[���b�J�Y��ɇY��w����j	�ܪ%.	�\�|��1�rU=[��!.��L�n�V�'O�U~F����1� z�Lohol��4m�ݔ<���ѡ���KA9���h�h��nn�3��Gl���H�"�� 6��� ��B	<���h�4�Ý��7�&�UN=J�T=="���;y\����:.�ٝ�
z��<���p���4s�p�n�}$F�KZ��{4uA��U����]�ڼ�&�ؤ��Bp��q^�`I>9����?1��
�+�sFK��Aӏ�~�iP1(��a\�;�{�?�0��O�'����y����Cz�x¶��%�礀4C�Wh0��^ J�E=2�y�#�垅f$:�=*C�o��o���F���:��u�TT]�М��ǹ�/#�*)��k�-�/� �Xr�D��p���Eo��Y�<����?B��Ñ��������:���R촀^�i��;�j2\�	Sh���HN�uKD|��+��^QQ�'�'��<c��Ăw}��	���2�]�ӄ�h���T�F����
[���S�=�_���U.j��H�&�?�g?�(��]�*S�=�������ζ_J޼.S�c�*u����Xc�TTRA�����^=�����$E!�
���{(\�f��=n8�o�F�����&�ȶy̛q�����6q��O/(*6�Y�:������̫qlR�Wz�x�qyV��p��I�Ľ
��A�t���#TV'�3I�_C���U�,wÀƍ J���o|�0��lK�D']S��̦�YVe�Š���7�/�ʴ�)-�C/�陸Su����md�>���>0�l��O;C�
�Z	�QG7_�@��Vj�'�Dce��I˨��M�rQ2��c���qO~���^��J��(���3�TT��pLq���^����n=��;��h h�mQP�K�	�Ax=��6���G>|�I�3���Ɣ���^�S�F�<���46�G���|�%�o]�s���3 
��| �Lr��L�-z��>&����_B�ۗ�  C��ک��Ϊ�0��EL�)�.���Ɉ-.C�-�i�@F':����ƨ�$� � ��J���ZV/�\Գ���_����s�2��ˏ�p̍�8���+p�����а��X�m9_�%�o\|<���Avv6?/o��G�3}]:�������+h���u-廴�]��{�������rtKV��c��7nD̺{a7�]D���,,���Bm��g�3��v6�i�ж�e1BREE\����{C�n����yy'�3��C"�����6��
	i���989�K�ZX�H�����"���m�h��B^��y�RMEE�߿NOO��a0+'羒����{0x���W�~��&��B���J��aHxv�!��i�"���v�%�4hgoR���	�w�u�l�%�/1-p�Gy���u�o��P���d�>׾1�a�^�����N�My����:RdV��Ξ�JG����_:����.��Ǜ�3
в���L�@�q;��U�Ik��ư+d����� ��B���WĞt_����6�h��I2��yOy~�7۴޿�;i�s~�3���u��]�	U���9k������;S]��g�~r�L�������Zn��<3���5=����v��Y��"�6�=�JLY}z��sc�����S,7��egn?3��Ԓ'{^
��/0&p�o���8����9gPFE�skm��LJ��Ȉ������Gk����wWrRд\e�a�>^Ȃ�G��t�x�I�`;�s֔\ԑ����c��TW������}�9���З��^;���f��}'b-f���<X��-��x�ga#+kxo%!I�9�֭[�`	��W��|{}e�!�����q�֏`cOmuuLv�%|�K�P�e1��HVI-�*����=o �o������Y3�U+��=@4��$����8JA�0�*�+�����2�A�S<�se���/����9|�������_���%V���"_=n8���Y�l�]�V����h^���I�yH���IMM�f���fE�����g3�9z��$��_��uH�.��A�:���b�w�DӪOQ�Q��}�r�ܧR���sb=�d��S�,N�,��&ưȩ4�40�ȝ�������=2i�0X&S�e�Z���D=�������G/�����n͗�����,��n��Ó�  ��|��)�[��x.*�7�~�b��%P��#F��`�⛚��w��������a��	���FEٕoא+mS^2�D���"Bq�V�핐��X��e}!��Ut���,t��6#�o"���~0v��$�]r[��^:��٪�~�U�);�՛�u�"����rW�,�zՅ�q-n ��5NQ���q�f)�LN>�]����
��|��!k�-��x�툵���Ǵƨ�*:,�Ý5[��.�͗B�ġ�w#.�MÕPCg��NS�����,�uQ�7��������� �4;����޵��h03^ �F���ڷ3FF�s�v�=1���i�S=�J�I3I���MY4`��"���u����~���d�F<���U ����p�1��))$0�jƖ���B���l�"e���#�}�ݗ���/�e��`�C?<n��>�l>�'&�=�����V��8�&��/ls��N���ަ�#bb��IH���R�o}>����:����~�����hJ�=)&`�_=�2�Of�v\V�����%� H=�l�8�*���<!�#&�^�X��<Z}@����K~u�\`r|kJVJ:S3O�zq���V���30T�Y ����gsF\�l;�e�
U_�������Sj�^�E4���ʯ�Į@������3�n�е��-s�1B�Q�D�N�������=Yʒ���Tq�Esy����uY_O4Gbjf�
�k�F�I���jA>T�H�*B9F˱w((脠e݃%�f��R���m��]��5��9d��g��0@xE�(�*��a���Q̟�݋��2_�j�{��q�e���A��_^�O�@����f� n���L-�ߺ��͍������������B�g^�Fb�n��V���\�P���]���I"�T�BD�-���ݕvA���}c{��>�	z��!w�䓯AtC�H�.J[��e#'c�/01�كygR�Ӯk�|�H�m$r@D-�MM��ӳEU�^�()�@S���;���L�؇d���
��%k�Q@��i�n��:�����#���ϔ����b��� Ҩj�]��������!@��ghɱ�j5dy
�?(�'9�_&T��H\_׊ʼ��9� �����Iu�,:uޞ��K~�\?G�gw{U3nx_�Hر'�����7�  �ND�L.��X� @W_�%����Q��$b|Q�p}����ݒ�u�P�/_?���/�t����qQ���ٜ��S9�� ��뾅��@&����O����S)�E�q�x7?P�<�CAӉ�h��ۤ$�mUUU����!�6	����׷V�a����'\^��fw�_3dH�����,f:)[cf_1Y�T�J�y��=5�ϝ���x,P����;�q��-A�v���OiZ(�}m(\���RݪV�����7������ogw>���/�4�4\�z0n��� ���4P�Zh�R]迂r1$9�<Fuf%w&o73�2�a||O��V�,m��ddmk|Pن�V�} �G��� ���(:I\]\\�����3���� $7h�z�b�'+�9w]�秣�o�� ��e_x>W�Nb ~�$bd�N�ɟ؞J  \Mc��b$t�6\�8��n���\� �)@k�'ZN ����V��E��e�b�\��
���!!Uv��+m���l��Q�@���;��6��2�����7
��.>kpf2L��%��:��U��~�J R)�)\5��������?*~8��DFcs����'�Τ��}q⸴�d�t��V�=��M�L�V��r����n�� �rp�--��v�2�h.��u��r[ �*ㆣ}��Y䍩��}/���Co){N��R�R���/��g����~gV!셥|�z.�T��=>��Q@�z�B PD��up������9G���1��#���K�r��H�o��қE�%en��M(@ͱ�*m�%���l�Ѝ�������k������d��ͬ΂U�z���K�+���OSM-LKv݀����R'�ƴ79�^n��6�uA�[̯�T?,�<c~���C[�x�+��X���V�NG!�tI]q]��1V�E�w)���,)� �\����m�Sss^����4'�ϓ�s/���R����H&�5���9�s�{PP�T��`�+�'��ʔFR���| �YݱSj�tr/��;'/��=R~£�e�*] �U���w!us�5�)QG���������RO�8��Y�e�>^1��6!��5s��LZgh�F�^��tU�����;Δ3�M��]�|7;[i�1�p������EL @sc���Z�'�	��~zѰ��>�LǊ�L7������f^��f*�s�+������&</��*O5�=X'7K��zv��_����X���1�ݱ�v&8�� 6�����b�i~m+Ȏ��	R�A��2pp��mB��d��݀�w��7�n���+2��5�K��h�L��zuoH  �� $.����@;�;Ha���G�2_6����駓�/���3q�;���n��������:���hbnm~�Mε~�6�f���'#;�����]�qqs��"�h�����=<Z)��(�w��Y����cae}Q����������J#��N-��8޽�,R���_��v��v Y3� �Cd��Bq2��ܯ�di"E�	�w-�+���|�/%��9{r0�u��� 2�]���3�}�<f[��'�5�0xئ��q]###��
�����* ��~a�0zqcK��cY�����<#��� ��]��dt���	O�x��������/p��Ї�B.�AԜ�:��]�CBkp������e.��̒���}������Į)����Z�i
�y�.y�B_&/(� �t�-��شr�a	
�+))]Ѡ��H����W�!R�"�<r4��}��*���ʝ�t�6+I_�p��V^���\[����ﳑ��Lw t:{��S=�޴��k� �nqqq�4�Fr fF�iY|@'K&˹���k���x$W�ƱRI8}X�'���-�+�@�ef����ƾVj=�bIE_�����Nof�����K
T��r۲?|��a���*?ڋ���Y�񯿟���&�{�ei�V�2
ǣ�ɖ癘(�I آJ$qP���]�����fŖ�ǭ�0�7~���S�����w�}&c��W�>��O�����c1β]q��zx�+�`����{�^m{ܾ)��~J�����:_B[24hK�4ճ�߽~	s�����S�P�I���%�����P�Bh���X��)?`x+�YK֗F�響�ܔ�<��m��`���I_Da�u�0��	@u&��䁍@?Q9=Z��Pu��dy��������"�O�h	5$��I&Hnj��t��鿸�,P7%�1�Yq%TT���?��+����nX���g�±�e䌯3�����'��l��+g�-�%9�]�ï' �X3:ݩ+0}ţ���Dq�Y�R��#6���Z�t@~�iu�.R�Yo��cc�
b��AH*���" �t��t,�t���4��,�)�  �,����������<�^�#�}��9s��:�̬{��9!C��Kh�^�5�~���t�iy�%El$����}���Ra��[	8������k�P���2PF�q�=P8aR�.d��SRQ�ȉ<�~�VX9r�^�MO~��(ͨJ;�~�OW��H�B�v*�� ���Vڊ��+��~ś��_{>@3��.QWP �3�D�L�5Ͽd���FR"|])���z��3g���a�I���$���lP�.�~�d'"���e�9�����>oߞ�9p��DF��S۟٪���[9�cވ�ϥoNd����3�&�$�7�'JX����KSc�%w�/��^  x�7r��rݶj1����RK��tvvv0�!
�
S`1P(7Xl�$/�g�öt���'��a:�}�yˣ�",�l�T;#�aa��9}��
�-��h�]�}��aG�B�J\�x&�ſ<������er���{�8��%�[��$���`�+����9�/,w'
�k9�`�����{OIG���?�^Z��t��yҙ�\Nm�e'S���E	��y?�6]�d�w�-��GQߦ \\&�؀�����L�䚪z�Ȝ}���Ib�T�3h 2 SK�S��u �eF�����M�^�h�����"9�'�$<�cSA�L�0��ߐ�[-�k�@v�$��Ԓ�4�]���'�4&�����m�T��E�Ԥ7;6u')�^t���c3��O}$з4���u�� �#uj�q#UP2 �[ZzzC�ut�������+TΜ9�^�^e�4@�NLz���cxfl��ы[���?g-!�vl��D�&���>�_��(ණ�a$L�>�Z=�r��
ݛ6_\����l	���oZ7R���7ByH�pEI�V2���
�eu��!H zP`�<Ľ��ςp�.%%�&X�*g�����J��['�/>(����G��i�d2����^�]� �\��,��0Չ��z���I�꒧��N��(*)�f��u
Nǩ`�����G�{�0��&|}?���ßZP�:qq��I�* ��h��f����kY�@uV	/��=n���MG�C��a������;���j�/ba@%0���H�T:B��3���"''�ܺ+F�) � `!�?���6���l�_߼�"۬�{s�ɈIn�y'v(W3z��ŋ@B���������W�.}_QML��3;F`t��K�Hev�o��Q�^�}��/�x�����+��`ھ����- �kX���b_d�	#�]����А��g�$�U ����}�"�ϡǢd8�T�ig�!,,*
�aY&b�V�\���+�t'�Bur�]m��ҷ	�}?��KV��6��LN�%4L}�C�ޟ�6|��Ý?���]t���w�`OX�ss;�i�nݺ�f�B�,��8@\M3�(������O3���p��J��ˮX����O�z�(/ �j1������wG�!O�~�+k������Fh���c���Z�*=0Xc�P_2=Pq�ߩ�@�I���f6�%s����a�4�!b&�e+�R����Ȍ�>UN.��(IIv����(�=(�S��k�&�� c �p�9����bD��0�MK	
�V�O�"�v���(WD�i��	ȷ΍��ͫ�|���k��P�����ǥÖ߿�w��mE�k����֕��+�W���+8mg~�ߝ�mWZ�A#��JZfן@�w�л¬�oM��a'�|4�hY<4|G��U�^�Q_L�5�7J�Rd�:k��v��N���S��OB,��^�qc�����2�|e��d�/���՘��J+4Y��-t�,�~F�9O�]�h�'����=��Ջ�j������壍K���&z��ΟD�gإ�bB���t�ߜ�%�+Ӝ�O��;[$�5�U���;:^��Hd���i��P�@_
�@+��:�#!)����ߞy�{c#����8�z�2�CtqJ_._`�uvb���1���J'�l����T��h��H�5��C������
*i1��G>�Ij)Ht���u��v��Q�BpZATS�y��2ޙ�f�%,��U>ni�d�S݅TB�������rZ�8��P�5��q�U(��'؏s��S4��P�\1xZ���5����0cw-�qz��~���fʀ�8k	�8�k��=eɟ޺��#i���2V�q\@O��S]��U���\!c���AHFxz��3?��΢!�U���b}��wg��~�Ў݅&��"3�-��f��nh*  ѡ!��\��]$P�SI�i���<�����8W�5�2�_�\�h��C��x������;�+y�sa)������R����+�,��l����[�J�A���U�H֒��Q��N���~T��;�-�V��G�{a11C)��^'���׬�&PO�KrM�q!Q�xp���������~ѱ�������|q탦����F�!�a�����'�3Ƹ��斖��x >�`�
M��+��$U4�Ed�}K�]�0Z(dAF�����c��e�O���6�N��g h,�7E�RX�]�Sɠ��kx�%V���K���ʵ����O:o��@V��/��C&�F�g���g�|�<�d����3�5��lv(�q�<�ۆ]���`��X���>s�,��uu�%�`�B��v�g�խ"R޿?��WJ�PY�[OO�\��N�]m�����{s��>ù�.%��1�����ұR9?~���������c����/x�YO}�Lfy��e����䯆y>���[Ho���&"�?�B!RqO�Ľ���f��H���ii�������>�O����r�>���v�n���I�s�rt��4�y�QO�=\Y	�y���N;������@h��Ŭ5����S�Ε��.�i?�^U�J�A��T���� ��۳)$)''��{��-��ˤ��|����2@�c%Vug���x0��#��Ā�q.Z(L�>;��xf�ʀ�Pcm0�a	=�PR�BT�A�@��b\H�8�����Q6$. ��ߔ8f��U�D�c
����Bw:��8�{+59Ef����C<��]�lnܱ�AG�w_�
E%��?����]ۭ����
]�O?��V��J:z�Fy��/Q6������H���<�X�\G"]<�>޵��5��� ���,�ʓ��8t��LB{���p�7_��u�2W�q-�T�Ş�x��ǵ�Bb�䀵f���938%=�Y"��pG���]#<=e�����7;�2>y�����²v�
n&]��*��\�, �����.�TV��+�!$ t��Q�����GyZ��r�lj§�~��~}�I�+��nЩsĪ���a!��S��P
����8&g��������U�a
��]��@K�ڃ��eEDDBz�b*�֙Ɇ�]��JB�;1V=Jg�p~�Tw;L!�Um�{�Nq1�R�c�8��ՙ`L�q֑́�wҸ��Y",,LMS���p(4"":��t���qjk֮���I\����}�X������m�А���Xߥ��	��%�����Eq�
��f�{������y�>�;�Z�}�P��-cU펮"���{������+�9�rrA@K8WkU��:�B y����(����;�<�r�/�����[8?T1�4xF����;ﳮ��/fpY�͛�T�a��_<*��4#a9��b�h��KNA�Lk4K���d����;L�mk���J�Ll�BR�J��!�����<� ������_�tU��Dۏ�[ȴ�� ����g��vmIuAny,=ÿ>�[X�$ ��X�"�q靿�A6OdG"v˨���؉'�o>=�ZfN0K�l"�w���_ߜ"�qc��Z#%���sMMM�؉8@��^c�A�}��a	����Wxo��X���y���F?O�嚘2�<u�� ������iL�C,�Pi,~��E%Mͬ�?�0fIec�w�60�����+�f4l%���}���;�x�>* �X42##��iixD֍!tx=mf~~�/r>5�"��wk�h���ы5&rkVAϗS�U��j��$k��J���H�i��*Q���Ǥ�ݽ�6	k�+-!..�@�gư��=?b\�Hh�0@�M1i0�C�m4�)$���u���fyw�j�Iֱ�uB��T���YYR��}?HD�@ �gHII-$  }O
��H=��{_��T m�'�ӓ���dG2y����;M��u3�ޙ��\�
����� ~5���4640rs�Dh��O��kN�f�e���Դ4oc�B����hz�Z���[\��*�~��	ķwU��_Vo�rp�m�,�O%���-��-FKV'�~
�ig���w��m_ ����
�����|�`h��s��Հv �{n��]����#��l8zm��r&�J���5����bb̝.�}oPw���!�=Y�bm�>�=��9=�OS"����^���;�s�A�����D�¡a`�Z����b��^�����k^Ȧf�O����aD2%}�I�Ym�yڪ��A��uE��ӌJ,�H�yj��S�A��ѱ��gΜ	�Q��g^�M!Zr�x� f^j�{�
pA�N��K�cv�^�y�ӎ=;�ݽ�GE�+l�۞2���������X��*#}d�u�f�#ݷӈ��Ys���%��]h�uP�֎��b����v{?�}�//Y��|��@�
�����[�op�|u�p�A�˾]�`��K�W�=��(�gw�ܴ�s\���E�T2t�G���|g�M�ruq=��TN�F]��a�u�� �������1c���(:n���(d���:y߽f~gy��ۄ�ⵁ�Z��݇��_�w7��AG`��y�jٺ���=�z��� D	zT�rW8�2���)$u��%}d��������%�@V�������}��=���R1��K����T;��
��0d������K"���m�J$A]���ɚ���y'ªЇ�rRA�^K��f�c�̖%���){�M�Y��Eմ�j�Q�}���2�""3_������m���v�Y�s�����ο����:F�Bf���˟X�yS��'�!���-j�/��|�UA�=;HxO�2�\;}M��$$W���A8�L�>�[Y��U�{~�̞���A@�K"�H��|�k�����14�3Rt�[!n3�[0��3���4>�'��6<�����W
}0S`D�0���l��A ϱm�}�D�A��PB����l���u
<���%m�9�����6��Z�����5�SL۔�V�Yd�HM�C-~��y�ٶX��ލ-�du:G�R*��T��H駉�e���u���TT�2d���?
��Ir�t	D��t���^d�O�מ\q^@�e����pj�#� pE�H#��(e��އ�Y�{h�2y�sD�׮�S�-�������?�����}CJ~;�D�&�y/$��^i
��Vr�cat���Nh�z���������y.��d�u		))��ҡ{�<Y,��p��悔YO� ���g��~�l(q�Xo�F�$%=gR�z�9��V�9!�����*0]����S�T�j5,�=I��l
�o3�\�{��x~���ڣ0�]��o#=�����<gu6�� q���n� ���P����V5O��W/T��?FkWX�Fh�5��Ci"�^����涶���7f����Pi����ga��[3>((��ۓ���fx�.<��wҋw��2��}����ӸD��r�������?�J����.�bhh�S�9`f���<uвV�G�!�����{a/��	�-��������|�kڕ�;�{Y`�+��Z�@������;�WJ�'>���ꗺ7��xoS�W���P��֣e&;��p����hh�o;Ґ��͹���`dY�D������g�\8 }	�i@�j���7t�f�=����G��?�ED�>�����^�+)6MYل���fz���0��2��h��B2mHLT7`�é�к]��J��_!O<A@w�E3�� :���t�T�h[!Ԭ~����>��_�&�w�Qc�y+��}��_�`�yWi�ܒ�Kga��{u��x,M���k���D��Z!]�|1�EJjCj����H��@����b�MŰ����1�K��V�Q���t����:q�q����Z�ɓ@�6��y>XX�����9q��{���A�6���i�KY�%�ƌ�Az���U�3(�w@�2;\Ѱ�gT����LI�������uO��F��� ubTN�3qe����}y6<��q��y:�� �99U(9����� �f�s"-����,+�����Q��*����G�f݊+xg<xQ��J�Ӎg��)BvN���C�����~苯��"����g��̼W����R8:� �����瞲`4t(��5	II�ػ�8 �cڢ���۞�f � %_ >AJBx,���`I�\F`'�}M�:��'|䩖M�7.9)i�'{�\�Y���n"�������r�϶����H��*�;K$��X�������|ܛB�i����$�S�9��0.^�v0I��s���O���dE!.}�b�f�e����L�����X�߿/��r�9:ޓ������N�*�Ff9���G�X'���-�r��Gs�@^��uuR7��Ǘ� ����>��t
��S���Z�8�]a �����⍂ܣ&��ȵ0)⤰h.�F1m�j�t�Nv��,�!P�}�������P�B^ю�牔T_�ǲ�������4t^=���ցu�PO���#�w���2&e ��Lz��J?/ Q��66��[M?~t��RӢ�n?IruS��r�7+��O��v�r��7!�aQ�P����r�� ch�z
��I�L�}�E�fu�	&-J����u�Z��9��ys1���Csmm��|ٟ{:v�)��˕��)O\y���]��ə���s��b%��Ӯ$/�h9��� %;��5|��<2%W�VD��G���x=op,���n�`��ޤ�w��{r��3gՠO�w�3�'���\]+�x&?�19:���^���o�\,���_�޶c��발u���1`z~����(�{���2�l�2)�bDD�[(
�����./!jVFv߿O�UⰢ]�3���%##+�[���o�6?y5+��yȷR���B�'��} �M6��g��X�m.��h�!���gN¿\���	OoV��.$!�(��T���
�T�����Mi+�-���[��JyD�g6YkWd=`���NS?I��/���.���n��q�y��o�<��g+p�!Rcy�૸c��C�?:�@IIiB*ɠ#-=NU�݊�g��?
�'E���`��̪9��t��^hxx�t,o�F�%``1F�ow OȨ�|���B�BQ�6Jn�N^>X�}Ǡ5^P�&Q�Ǵ^`��`��&��br{zEeeܛsT�{�7���
is��f��"�H�Gaj�����f��#��8�'^ v��Ы��8�j������+~���G�z��~������6�͗(Ҧdr�̨l�:��1��k!������0|�w�����y�\NA��U���6~&._����# ܺ�~�Π�_HV�}#����X`��AtZo9�r|��ʪ,'�{EEq�O�_�xO�m�r~�>pMX�g>���,w-[�Y���T��^�/�4�T� ���c	�˟��w �~����c��q�� d���Pآ"6��E�Qm([�������W�
ԣ��
�*37w�}o�Y�4t���vFww����b^��.b�'[����[⨦�O�>;
�L�ȍ=}�`���фY�f|�8z��ıxu���-C!�&$9 ��ex"��T�Q/%���K2,LI�󱈗I��+TAq�gC��F�a�Դ��Q���7�E3���}
(>>~Zd��c=��eW,wUm�� �ʿh_������i���o�5��}v��q�H]Ͳuk��X^D��¦�h�|wG�0Ԅ���ji�F��e*Ek�< ����B����9�zo;
�
���WH�u7��?�����/փ����%��^�s9b�y�%��bdsKU����"Sl3=�k%��݉�q�P@��o-������\��o8���^J�e'�@4�9�}����r}�m\aq�ݪ�Y�r$p(l�Y��\FQP��{z�kU��Z�� V��f����Q	k��i:3/)������֠%�9��Y<v��h`��3�$��2w�6P�Wyst]�tj�QIQ;U�kz7/���E�"�����:'���ڴcP����
M{�gu���7��&�O�z�rۦm�!Wl1h�g�}�nx�!>ǣi�F�2U{������Qvd�M<P�=}K�E���@[m��3���N
��r�-��,��<�"��v&���>�QJ�a�v�ٱ>ٿ��3S�"��|E��}f��F+��1J����ꖍh8�m�#��;d�x�`V��ϓ�o�={�����������U|�n)�%���=�����r;�|���=��܄Yvb����k4#��������B�����p�l�`8�1�3��R��dfeuk9�B]�n{�E�mph�[��C�#���U��k�P����� w���A���H�z���x�����i�+���82�X��{/<[�k�䊪���^��AL���[Bl�zX<c<���Js��l�%W>�I�,�����Y��TXcV�2Sq�c/�Ta�ꏗ��8�X���馄k@!>�.�4��aV���K9�ژ����4�J�3w�u&�X����A�	�m~8�q�uV#�>�W�Ng@@8=;�A9}#55*[��򇈥0��"����,����h%;s��<����l0~�+:Mkd=b~�P*o�.��(Ry�M�Z{Tl����?���A�wjy�{���Vb��F��g8�?"(È��qjĝ�����3�wF(�c�L'���/dW�M�����v�,����j
QRW7U 3�ߝKv��D?����b���ӓ!����F��2tf#�t��c�mUZ�rѢ��%_El]�^���A�D�(�����y�mԅ~��E�g/����*�Xk�n(��`���WaD	����٥�t0��g��iՠj�W��+��@��sEfs�Q`�121�6�A'�ܶ�әr*��@�y�;��9d�R�ØTv�V ��3�������tvPAee�Ƶks_��:������]7�uB��ļM{8��d�a�(M1��">�m���N�%�Y���f�e,�nN�ڹ�(�9�	����x��
��T��'�W���U��<�Յh:�j�-��x^<��.�s�tg*@��eU{FBF��Y��pf�$�3^@����^��� b��sw�g�Nݺӈ�������x*�t�+5myR�S̯�N��WZx���̽���y�C�̱�ǧ�2� �]�����1_NfY6DEZ�����/Ə������n��R�~�0�����J��e-�R��[G�z�噳E�~]���k+�n�qYw�N{�x廡]e7<z���r�0�V���s��rrr��u���'��(�&��~����������Eq���e���CGM�c�22`��+���,i����fo8�z��@�4��ొyyyj���P�2:	��0�uǧ�V��Y5366� �%�C��,Z�干�Z&p��:/�B���*h�8ԛ�`���?b���Hf�w���Iga�1\;3��D�����D]X��T��F$��m�it
�n��Q�r��򯹜���{�H�	���MfLdw�^	e�g��,f��uF�h�&�ߴ*e�.�d�;iY�qL^�,�	��ʇ?��;���.&��
���6���i�e�m!j��7���gBg��: �"��:Kw��E//�>�k�����d�-v��6�6jU�c����~d��i�*���P�|K��Na(��l"'�sE������xB�8R�˂ ;��r�?����8����Ž�݈�~?B]�������(��O�l����2�JgtZ�J9��Sv1��ĸ�?o��q�쩖��-TP���S�.�ﮁ��'��G���"18
�]����1e���E�ů�&L������S3����{��o�E_#K��!K��+Cͼt�; CDak?�Q���	���y�L�B�e�T��Yom�/���mPƉ -�N�3�������v�3[����(q��y�{��]##�����J���T2��?�#�>��F#�¦!�~�����#q��?~� +!�t��������B��QCC�Pp�ڿ�*:� �����hPW��#r:�V����R�Ą ���ze�cg�L �8r�E�?zp]���M$�p}��n^��1U���ì)��5_��	#�S^J��-���cqz1�ȋ+�Dp�Ա�W�g�S��'%=0��=5�#k��b��PA���緭���כU6$�H1�p�"�#��$����a,��>�-��]-�����qv���3,44#%��%�����*Vz yB��Y���I��ٔǥ�11��$���?B��ӛsX2Ν�%��_nH�?�")�^����K�;}��h2D�V��ͫlt�˰p�'��%��JK?[S��D%}z#����NZ 7�<ؒl�Eݱ�3az���\�ӝ�E|%/�nDF�����Zւ#.�<��o9�D������>�!$��)�-$���:�����A�m��p̆+� pl.1f�Q��Ѳj:�cj�^sbP��m-_��d���c���I�UO� ����� �O����;�Q�Q�7�a�����Oi�i	j��݅C5��b�e��^�B6�������/���K�ڇ�"�J�8�b|Z���!
؟GD�	�����l]*�-�򮤮�$�\E0X���~`��c�3�5E���Q��FF��[�A�go������;x��mvy��0��ʂ��;v��NB�rf�Rf1�O�^7a�ݻa��0Lㆢb��D#�UN�F���5L���d�2�"qS�T%ϷT�kj�q[f-nr?��FA��dD�\�W{޺�񚻟HZ$�j<�2�@�2�w�u�p,�õlXv�`8����{�'��A⨼cW|�3�P�m�"�����KiW|8�bm�4P�F>�P�-��5���^w0�܄��w�$�����Te��~��O�R��e+z8B�B+�m�\�)|�����Ȫl8�a�gs�fP�u�2�#�H/�҈����K�Υ�Q���zd�I��lO�E(�����A1��'|�|ES�?��Y�|f	������ʁ�@�fy5���[�m&[��s��M-��S�OY��
���� �Y�/!2_�X���_1r�+����hK�P?޳�9����]�u����.���E�O�^ 
�e���K�{��:���I��f��ajަ����o)�C(ڪ�Z�O��7���壋��+1��nCŹY�D�_�W�}l_U��+a��C�w�?'%=I��̦��FG��"8�4,&y	��]�%[�*���U7�-7*��Yv��`d�L���q����tHy;�"����"�.룳����y��*AN������=m��c{�$�>��]D+h��ƾkM�%��)M����']�/x�8P0H�p�1�#��V�ˎ��ԧ��}�>4�����f,W�+� ��=�_q���"��>�[�a��:=d�2�VR�q�-�z����F	��߶����Ҳy3j�j"w!I!j�n�L�9��√X��T�~�Ǘ�N�s��s=��G<���+��K[��d��s�Y�]��\�r��:.�	������8��:J��Ѿ֓�v@�HI���׌�8���Xs�X׳�:j_�{����ӌ9pSB*OϱB�����S0f����n(t����$;=�ɴ��������5�6.v.E��o �+jJ�������<o�b�Qh�.�uH���2j�A>B\F]���<QWW���_B��_��֐VҮ�!��a��f��fֹ#r$��w���G�hes��$%��8~�����?�1[��_g����<���K�$��ݳv�����&oS#8�+�(���i�9�w!k|����7츞\EN�9�[���M]J���V�J��Fu:��~��濛/��!�3�{ϑ薇����4����&u{�:�/���糸��X��3� �z�vS�"ch)��o�v���	�|�ʆ4���|����c]�I)�]f]>ї�\��J��KC��悚��.�<!!/*��������~��_d"t֊j Gj�3�N�l[�������D�	��f��߇�[����*���2��l�Wod��|gM�9W��<y���3����M�dm�-$D(�rϸ`s:����%j������[�؞'�\E��tՉŬ�͗1=%�U.�'��t�?�S����T�y�O�\a+)%}J���a���$��ܥFr�҆�v`�v�~�;�:md�}_a������������c�бI���4h����
��>/>��(���H�kW�TD�>��<���|AXUTx�v�����	���t��u �w28}����z��_�Վ+��cE�Ra��"��qG?�!o�^}�Y����/��Jv��Ӑ���x
��f��j�N$P�n8��zn��ϝa��}�W�;��!!c[ͨ��{��,	�{G7������pa/��>�a�ʷ�	�#�ȯ��;�엲��"�ll��Mca$�)!�kF9)�����>�fv�F;�khx0wM=,�����x?Yr������JEڹ�&V��]4����������4�c;���׎�R�y��%J���u��.-��]� 5�k���ڵ�;F����8����K=O����2 ��������<���!�c��^>L��Qํ��z��(}������*+�ه�/])r\�8��^|�RƯ��%>g�L��t�mt_�����˧�KW'r����ѕ�sZ���������d���wg`��͙0ܑ�Έ,�����O�4ٴ�Sm�N�b�u]�YnE3Lc���X	����ʪ�����:����"-2�8���t���zE�E��9��Zih��Rt��43�?�6 ����s��;Ǫ������H��Cޙ���{e��~]�k�'z�ϟ/�ڮ{��?-�V���;�;<ꚙ�@��Q�����u?��_��y�D21�Û�Y~Е�x���cu���:����uh���#���۴�p�r=����~�C���.a)��Y޵Nrs��ɞ�����c�����]��n�]��K��)Q��ق�\q]�� �i�3�%k���8���aWn!+�$BHk?@|��JK^��h�^���Jì�,Hc��/�+NAQ�&���Ƈ�o��_��4X���pZi�gk/��Ë����tp7�L��g�Q�N��G���%	�*/��3*��t�)F4rr,y�]�2
��$�=%6n�D0Ō�.֞V䖙��ۊ�q�=y79��5�����A�ϥr�v@�h	�ax�6�0cՀĉV���.hc��XF�f���q����OJ���:u�a���C�/CT�%�������#ʆxe_-�Xx�jmR�-t�$=�}��?��f*L8K�A P�ALFnj��yO�fl�� d���厾Y3u�2��@�E�,8s�VQ��_n"�V��N������HY��Q�W|�g#���_$�`Dv/7Ɵ�E�:9���&qY��ޚ�T֒�]���*$�ۇm8��rPo�(��<��B�VI�~�o,���:	�9.-u�Q���-���G{�IH����sj���ͳ��G��7A4��j8aKQ̯����s�x{��'$^���5C���QX�%��":�l���e�҃�ā ��Fߪ]�嵫�n�٥`-1X��N��GKk������>9V�6����2؋ʹ�%��pfc�:����8�����w��&����y�������)8��s���n������;61�߁{����fy��b�!�������v�#�0���q:�"���N�kԷLm�c���޸�K<z�+���0���w���~��?x��&���������u�2�f!%�n`�X����*��vgd��[��46�٪h�en��Q�ӽ��*�}~��?`��x������Ѩ�[Ȫ�PC	8�+QQ��fٱ��]J��+��ڎ_3J����%�#��}T�O�R9�7���gw#̕�y�2/�
���We�l�-�@�v�p9�Tg��>p'��ok��F|R��=)i����Ō5W��Mg͟>�Է��D��m��Ŭ����?�jG����T;���^LPm���r쐵��Y��:��{���
5��\��^`XWj�.��.L�����9UuN��^�i��^�p�oRRˌ��ր����$�P���Q���j�0}������6�K����NB�{`=N��7c�ɑZ�i�g�}�����st�Mt�o��BP96�?��+/�hi����VνKXQ�'�5"7l����LY
2%*��g%E�KXA;w#ĸ��QNʞQ���'�9�S���o�D�,���@��,T��f�k�1����J@0i�(b�����{�)�`Y���օ��^�B6Э�U֢�]0@�%&���u�[��5�z[ǂ/09�'X�-y4�N�5j���[�~��D,f�m�Be��L��J�Lt���Q�ۤ1�V�g��[����;�A��{�%�`��s�nɼ`r�BL@]J���A�T��Ҥb����̹� �	�O��%ݟ.Ss�i��3e��7�eZ}3MtKL�q��j��V���J-�9s���%SQ�L�=�`�YT�p{3����E+v�,D��:]�\�J}G쀏�,���W���wA0.��������
�Y��;~����x�˦cӥ��{+��6T���wkb��H��,��	�o^�+Ze��Y]f��;��O���1(%��Sj�_4�rP
�nB����a(�U�<����/�@e�B)�.?v�6Ĕ��ז����x�HImk�JW4���3��h�|��Ҋ��k��;�Ĺ�o�Vn$4&��ͦsw�E�w���+��^��az�p�/-zu����A�]@�oG� K����'jM����)CR��ܡ�{Z��n�"^�p���8�u�ͬ\�
,k�r~tm��SxloJ���R��馞im7L�x��Ș��K.��mK�?.:����!Rʙ�[&�ɇ�@��lի7���hŢc���q(L���S}ݥ�L�����:TN1tg�����.��U��D��%
r��s�QE
�D�O|��X�ɥ^�PGǼ�Se�ج���/G��X��}"�QՈ���6��iQ[�^�#�a:y%mfg�%���ف�\(�b�d�*-v-�k�Qz�}t]�=��#�"�AX��Ԁ�NӐk��U�:�rT��[����5�h�����qg/Qg��?�;A��/����j�����qhj(��ѩ��㼻5��@8�*��Y2�r��RHA^g`�QllF)�.�[��=�m/���-�,�B;��:*���a�d�6�z52��(�����7�-�ZLk�� �rH�8�-+�J^;Ǯ�r��L����~dZR��a[7�d�q�U���Y���n�l�5Ldb`j���L	I�!6,���5���[!)�
錬�˗�22v}�%���zZ�j��{_�e3�x��]��.5&(�##0�r��{)������)��,��g"��bn�!�-Q���5H���Qy�@�4x�e�R�B��*�D!�p�0��KU5��X9w��.�|>��A܃4�*Ǽ]"J��V�q���r��H�ti���9���f����L���3��~���G�}}}=��ݫ�7=W�͹�n>�N"`�^y[���*�fQ&�4���6iŽ��ȏ~txR>UN[�����Ft�O6��ē��Z6�Ǜw��W��f	0 ��.��3��Y��a��p�1A(������`*��>d����X�}|��׍k$䦈ې���S������ɑPA��T`g�T���p�|�u�T�U���=�Y'O�#ҀEqm|+��^# �贰� �y񨐤b��uT���:���:e���b+f�H-5�9�*zУ�P�:n��ˆ#+iD��f��K��.;0�.�S{�w�>#�;��'?*����ˎ�
��V�*t��F�0tm����k���&��4M&޽���qH'Ι��,]�1q�ػ�}T� �ͫ�j��	Q�x���Hm�R.5��k���d�FQ���|��<�>���h�w�jwO֘1W�s
�Ig<^� oٔo�2PtsO�&^�	�<}1h�8x�	��T4����#-�q��A����������Q�F`	����b��@������b��.�*+
���,�\���$��I͓�!X?�`�W*D��A'��Q�Z9��YO̿����`8���T��(��}ҋ����[F�K
NUڭ��&�O�~�;���MV~��턊����j���pYDA�ȡ��&@mzK�%%���HY{�s��`���lp�<F�~9�R$�{x�|�e�����'��]��9��ny���~��1Y�u�������RXz��j�o��^�P��&lyE]��>�D!����"���@&�C8�u����
���1Y�ʢ1�_����A���� ,2Ó'j,ꅲ���Ef/DD���{K�'�}�6��������q��@��WOA��M�E{�Jm���o��E*��rw~Ȇ!�+h8���U�n�Ssz��)�n�]Ē� @t�d��=p���,[�n΄��T�/�5�t�1@�/I&t�����Y�w4�}b9�/IG�PU`e��_��\���q�������Y��9ӡҵ��5���g�A8��ߧ�%8��Q�?;�I ��y}�;�ӻ���6���� 9g�M�� e��r� k�5��b��tP��ƅ�H0ϸ�;�_�dD�e,�Ӏu��*�����(v�FTIc�c�����,����0%K�\Cup�fkUc��/Kͳ�k�����iM���{`��CF���0������h/tLzl��E�%�>��oߞ�;�'}T��u_�s�Oꏡ;��t���,3�&۸�w/�t?3���b���{?k���V9�63\�^�:/����tI��$��,����ֽ?=���Rv	p93ĵU<�@_�/�� ��@P���:���ݻ�OW�� `s�}#�ݹ��.�}�i�� =�^��+'Ո�j����ּ�[X���q+��f {�o�,����B/���;~�L�k�7�U�p��o�>�~m؀�Ȫ1JE+�1ʀ|�����9������')�졽@M��;ޯ�{~�����`�T������h�������!�c���/Ϊ�n:O]0�]�|T�{R���s�"���P��[��Is��@�I�� ׀����o���q]�o�S��T�	[Y�ec�s]��v;�����d���0���-��T���x��u��F���{����nt�*-U�
l����������k����Z��_22*н�ר�X�m*�<���/�_A�t	�U��������U�߃�`Kb�*m�[����&����f�4_ٴ��IL����O�)ogWH����\,�J	<�e4x�z{����PU.���k]10E�A�� ��KA���@���.��H��r����o��w����]���13{?����~�N�og���\��˦�@�f_����Fjp){�$�iKG�@���%63RP[�E''���@_ߝ��5��� 9���n	����rF�}4t�0�����n0����P���5�*�R8���L����{r�H�I�:]�F�pX�8���K�y�{usYv�\�XE��7wy�f�\�K����S����V��l'����!<JF�����Y�Z�� �o.#�j�a��:���J�]''/(.f�������*j�7աF�P��xަ�֨CxH�Nf�l��Z�a��p�SQ~��ɒE�`o�4���T�|OFǙ���r+]({��͹w���/O��R�`^P�&�x*�۵s�P������c)åy��]�)JCK�S6Z�o�6�V2��q���IC�1��;j5�%��bUr��E���B)�/>�(M�#�w�R�Ҍ~|zQ��D�EFf@��\U�:U>����*�_u����F�+��2vpX|�R{jGк0\".=f��^;{��u>�K��JPq&��dčb#��m�|O[�Pp�Ҕ���^QI)"��I��Y�QX9�e��>Tv��,���LR��͊w��&�u�D���8.?�|�g9ǥ��Ҁu���h(��Î���m<kI�]R,��wޘWD�ݾ}�v�if�z���%�v�K�aG<�Ĝ�}��nS T,t��K�w�����d|j|[�P�ܴ?��ȫ+������ɵ.H��/�u�h�?i�jx���t\��-�������b��n�M���9�HԊn��������uaG?/:��v�(�0P����_���=�) ��_�Ǽ����=h���$s��'f�l� Q9�n,S�G��<Ixظf=V9��2��+ɧK�.�ՠ��44bɜgoAC��� ���?I�n�%��}4�1�$�Qc�n4�Y4������u���^}:��<]��)/"��#a3�=C��aO�s�۟��IA���4�D�.%�(���L�9�;gC���2���in��h ���I0k��ë._N�7����x��[m�	��m�6��7�)�k$�aU���,�Z���A�M��ű�9�'�^��l���֣�{��X�8y�矀��.G�H \!������&��%�o?�9��*ݩ���ڂHyddWW��*5�h��\�=I)�}����nA���t.X�ݭ:\��ׯ�MΞ=[�����$#���g�������+m���v�WP���y�N�J�(jc��1��WRP0���ඝ}kmcs�4Q��
��٤��A��[#6�W��[�i2D�(9�O՟&W��]?Ce,1�U�**T�I�ێ ���r�J���3�Z#M��k�y"V��ǡ.�?�N>}Q�s��,���a�	RS�t��Y��&ϖ�i������&�U�z����Ft��aU"�`���ʊ�s͔	a�V�o`��0�%3lcmͪ�t�msЀ����<�M_j�o�)�Gl:�~�A�$x�V���wp[�455�a�x �����	>�BQ{Y�Z��A{/��&��{ d���.1���E���]����Ll-��_�H+�Ԛ0�����f,---A�W���8~z$T���ux�_ �T�Ku![B�=��r�,**
���7�D���BktQO�:n��+�T}� ͽ3�_dԝ*
E��Y~��D��4K���%�a���%<,�U,,?s
��Ԣ���J��{*�nK3�O�:��P3(�>K�[[S�P�*@�BK^Eq�>$4�٫-�ѧ]UI�v��'�"��Ge�DDL���_@����s%���`ś���� ��[��fg�^~	B�te� ZQ_?j�Ay*g�_HP�RѬ��J��Ɖ����������t�9�-ͧwwD���-�z��`����7q6�c̻A�.�B	7�R?#�s�]��lM3HpS��������ϛ�pQ���7���M���cv�K4~��	2�������6�����JJ�G����.�ݤ�K��]x��gg�����mfK��Y��2����^����rB,ˌ��zA�6-�� �����_�<���\2��qE��L�MT� �C?��^��T�c�


���6�Y��K�x0叨��<���	��E]�al�$e��������"���Vz��W�+�(2S�*��,��Ϳ��̰����D����K��[��+�+Et33��Mᄄ���9��
�����?odZ0xeG%kk�͌'����]���pL{�a��I�E�8ېj-����qqy�9����ΤW�+�׃��ۢ�:�ۺ�rMq�޸�~q��SݢFq�F9W%	���R�gZq�#Q]�4	��RLŌ10� 4,E��ؕ�=rG$hV�n7��Y6`�$[���2���*3Q 1�A��1 ����M�~���u��������0N����!�LԚA�s��	�z m��2X���M=̠���Hu�:v���T�8N�Ee#}�J��l�[A%���j��$���!�VI�@^�>�-Y�8.H����WRJ���K��-��;~�B�QF�t9��=>\�Ѡ�JCBVXX��a�7�3;�WK��ʆ�b�+���;�E3뉽:;Zj��W�kvW�=4P�Rq�p���H^���,@ ��O�ulԺ�~#��mm�#ROjh�G�Y�W�q�Α�uL.��qv��A�����C���g�aI���{?I��]�AE+���B��	��񈕩��0�V�AEͱ{��� �gwf,�I���=�Xn ��>�C2�[�.We�xc�c-f����l�%�Ε/����� �|�r�W^�N�����c<,)�ڇ��1�f$nҹ��l�H�&qƚ����`�_:/���6(���l�s��B��el3����!!!X���;��^][c{��-���� he��y�.�V�5AA�k��-�O��.�H�����8>��R3���L��,MA���Ϣ;��l&���z{�s=9���M%aa�m�l�$����&A��fJ<�����i��^O 1&	�[��V��ȹ��"�fU�0���Y0�� v��Q��h���H�8H��N�~��$ ��u�� � T�<xd ǘ�9���^��\����'{fQ�B�k������TI���Q�#6�������V�s���XՔ��3,��G.m�Ti0��g߅��8�r�<���p\��;&�����z͙B�z�b��9��4���,Bk��Ȉ��C�HI��5�y�ﺽ�9����).���2m��qeu#���AW�xlg���)��&�i�v� ���@�Lsuu5��@�m��X�v����=�a>ݦ�;�tƷ�gB	��sJ��>�'��q�x�xk��o��a��hZ��IMM���g���Ƥ�F	"33s�6�(�y�:e��K�.�R�g�+�����>"�r@��9���˙��Zr�;���e���W��nҺ�&�6�6o�����rc���y�t[L����QJ��ظ�k�Ap=<�K�4���'�z)��q�,�K�k��_�:�%㸃�h�Wd1��%�Tv�|1��A��}��vV���S	�}g����x���ũфo�IN�t�?�j�w��9��� u�y�V0 E�gs
j�vk�@4U^
�����Z6�y6썐��b�\�onH��(w��xmS�X��IW�SU�- �`T���(�j� 8&�;�e���*�3��Fզ2$�,V�%E��β?Q��f;_����K>�MRG�L���y�5"�*���o�4>Y�QO:lf%1�j���+,��B)�\C����?�e�8ĕo���-��|��?�7��3��fb�QjfQ�44̿v3S�d�H=���>��#���P۵�9m~�`SM-ވuT7�>u�I��q$��]��2�f�H�����&R�9���(#��M� f�������Yę�<���R>J#��)r�'�_(�vE"�5�$IWD�m��*/�A�~Ri>粿Y������1
�V��A�/u=�5���9�xSч�g�[���[�	��63�v#(�
[T G�b���P]���ۮ��S+��W������;����Ԅ�����E���𰰰�o�+ܿ�J�������W-�1ϹOEW�*.�B�'��u�D�~z�+=x�����q0��{b�YYY�w�yY���_��X��HU��+)��JHӖSN�\�r�S�{-;���\I�~�y%�d!ܜʞ1�`@ zL։���^l%�kL:�c�Yσ5�}MnY5z�*���G__�;�ݻ�+L�]��8����Y��|l�/�S���.M�.Q�P�8��.<k387�
u�9q�	C�=X�cnd������ط���ːq��BQQ���eE���_���:̮��t�]��lu��(��?3���f�G���	>�SO����	�t>�R����Am[��K9W]�^��ư���[ۿ^x²,��}�cI��9)���,"��f˺����P�c���|yP��=�����t��	�w��e��*}��p+�}2����Y£_+*�|�SPxI��l��G���	|�jv���~��h����`Z�/K0�JI������J�����%</��r-��U��Yn�>�E" �������p����C�y�Me�lM.9B��c�1{�-{���vn��!I|�����݂��}�|э�M>�AC~�v 9��h��X��l�؍��^*rq�\�+��uHj=p�H���XMWTl�&�G!���g= �^}���@m+a���m�A�C���s)T�c��ǐ�;��rs��a��99�dk{�R9y��{� ��7f�Rd8�=�KPC �#�5/s��,���1��mM=����G��[�{<+iͬ�	����wzY�����Ge.#!�~�J�G:���2G
O�z��|=����|�u)�}fvvvSIo��y�L��� a��@�YH` Bvwwk�=�*H���tp�Q?����m���+a5��,���Yk�q	��V+��Ǆ.f��	>
�VR��>�P�8Y�CC���Y��Z#�Ѐ��G��Q���̑��Y�I2O�]W�N�i�@L�O�d�Z�"�{�n�������*�)�U��9���'?ζ[�x��c2����~QIL�
�/މ��j�s�H���D0j��Ć�NGp��LA���������rʴ��$�t�o���G�c�2��Dߵ-ܻ���_�����kw����{8��s�C�Z�b�d���ȗX�+�2�U����:��U@��xW�����$ָؕ�q��-��H�,�c57���˱L6���*����y�\kx&s|i �
6��Hkֻ3�G���g�K��ļ��wviӥ���o��N4l$��4�g��N��-��Xғ�*�?i����&,�N�u!}���y�A�c�Q���[��:a�;�2�s^7\�Fԛ���[;�n455!ɾ'�;�S�.$$�t��;3��p�	lV��/�f0�B������k�sۄ�5S���8�UAR�\@���t�7O�Lx
����L�A�,1C�v�!��o��> ���@��Y�d����2�c��x��C�~Կ�h�>(�糨�/mimE�=)!*S�(��3�7���`����n�����pw������.�n	ч���U�+�����8��b{?>&&'�7��_t8��a�$�3ye��ǔ~�'&&H`��Tփ@lwO��֨O>�����Bk;���ƈ�7�Z�{�gM��U`Z�a��r�gC��ˡ��E�3Q�P���j o�d�c��Q��HlA�ajN�C�S߸�:����[xܨ���;2����{����ƾ���J ����o�z��4y���j(w�@ɵ�O=a�:��O0k������x���S�T'���˿����K�#5�}A.��Z�/�:���<xػ���+�3�7/v
��C�����[#6�d�?�!��5��
�\��մ�'���
|{�£��LA���3���;�����L�CcAQ���.�伾R� +|�,�X�r���:퍋�I�nZ�C�d��D�)���ɟ�2���bpO�?�]�gſ��i� ',��Թ�� 2��o,���q�N�jK��8S� T+3���@+�v�WP%F=�@�)0��Gl^��/�ɤ�tWJ����n.-��<>.n�
�~t�؅"��	_J㦀k����g=vZ�	�	\���\L�4����A8�FV@@ ɀE�";�Pc��o����QW*�,�DR���L�vvյB5e�ƖLʣ488�� �P,�1�8u��l�AO�$�ƙ���9��Z�������������|]�?70��	��#��*n�(JųH����^=G���n
�+5�|F�)�|~;���|N�}li�h*JJ����)\����Y�ƽ��7�K<D#�����3�3�9��Q\��	���+�vKc�u���zl�-����_c~P'׊��G=�o�=��8�`��⣢���\��RJG�y��a�r�g5�D��<�p�cu��p���I��fC�N6����n�b�:VFL�+���O�5�b+�ѓ�@n}M>]�]��y�6��nB�hi��{��=����ۺ,�jaj;$lq���[��la��-�P�rT+�G�:��:KD�y��~{�b���2��_p���A�+2��=ٸ;�ع~�2>5�,F��Y&�v�F+����G'ܗ`w���Zթ��>�g���$z�6�>l�Y��������8 ��ww�)Qʻ;"��+#6pk9�]MV6	n�ö�(ײ�<8��/��rA�6^*Y��͋o�n���7��}{�d2��-"��1���-��C�F�	\~�;@�`gv�#��[P�ޠ#оjT<�M\1�c����/�'C��'hj��ammݛ&N�T��+iii����\�ߛP���Z4�9؍t�m���S�|��g-~�p�
nԀY�0�:����\��\�F�%g��"�A�0:�|'^2(_n�_�f�A�����z�ذ�[ �����S��ed�~3+�|�?����jO���H^�X�������������euyv�JJ�#��m���G{,�,���	)v��Cm<��O�Y3�����ϋ�M]===�v6�TZ��ja���RKMr0_�[���Ill�ZFn%�C���9�ëu����S����vj�����C���p	��5M����|���5OYsax�Qv{+H4X��T� �a����'��]���ź��Q!7���VC�Sj����Ѻ��1+�k�?��w��E���Q$�Oz�������wbk[��O����T�̰���d3+�l��e��1)�I������V[¨i��2P���5-�ꥦ]�͡&q_�b�|�E�m�kh.Q\��}(��K/�y#h{d}}�9|p���~��u�LlN�&¦ۙ�ɷ'��5c�W@~�u��j��n���窦�[��� X�^��q�	��&��#NۋE�}�_�t�-��Rz"�ϫ(Z�_�gXd�	f��+^�M	�.,�M���6�~lgg�ҁw�Ttߪo��0�Մ���+�=�"�g�I�ո��l��X�$g�|��\�DT�溹��qQ�����6mlCU
����'�>�f��j�����x����5�g�0�X�Z��@�H0Y`%����yZ5ƽ��I���phz
�A����%���eZ�(H�J�b`sv�=4w���S�ɜ���~��w�cs��a��o\��˂�v�@�wv��y�f�D���!l�徇"7�s#���[4��\���;���@��~����k	��7����}`�#��e�_5�u/3`�*6��p	 (�8EM�<��N�#|�Ԑ����tTT���Њ&����1�ȉ��r�2�97�Eoa^P �ϖ�j�\���e�	(��A��b6�����m)hi��2+	RMY*�y������<�W�"
�t8�:�9(sP0�n�7�y��R��iy�ہ(2wE�y�S����ᾯ��b�� ��Z7������Uk�뢰�����όﲗ��O�|`[X���m;{3�� `�!2�,�zM{A~~?��j@��W@f���8<��[nYB�(1TXX�۝��xP�Ɛ����P\#ȀTAQqD���䮉�C0`�L�e.[�.�%�x;7�k���p���063R�L7� �Cm��M���' ?n�K�a������J����\��Vg�!�>#�p��k�;`��hBZԦG㢅J��E���>��d�=��o�#ö���{�*~)�'E�����S�SO%��y}%&� j�����OMMq;.�(:x�������L HV���+A֬ B%��@F��pw����\�ŀAJ&E�s���#E�kk0��&�!+7W���q�֭
�0����w�< �b2�^(��~fa!3�Ƴ�:�M�����Ez�4�B	� KD���BL�7�6�<��X��L�yV/<����_��ݲ�<��Ld/�?���\��I����"da05�>�@�7�p؋��Z�q�@���~��:����}��Bݻ7.�$&
�<y2=��
�Oj*E�1qNy��I��_�n�@�3 ��:~��E�� 7����9)���%�^�笋�,8�<�KQ'Y�����M�E����C��� ��:1m>�(��p�lv�3��L��:*U�Yu6<̑�:�"@�N���Q�nM��������糹�S�cCZm�\�xr��iT�u#A�}�x�<x��G0q���v��e���x�E9�a���^!�;m��ߒ�W�y'��R?�EX� ;�A
x�?:R\]Xh���}%#m�i$c���[�'���ټV�-ޚ��c̡�c汓G��9#��!���N��	�����9�O��g�ARJ�X��#�$�H����]��]�i��I��v�ڵ2��Ω�	�i9�Ǳ��K�^x���.w)��]
�vJ鹯�	m	��j�pf�^ng�V����D����B��"������ᰝf�Usuj?̆��&���A8~�CE>oq�F{�z$��SA�Z�5�Z��3ka��uz^/�u�TK�S�uE2M'��g�E�� �y�s���:��9�.���
C�Bb�����?N�镱��E z��9��J��z-�����
BZ�� E���2B�MV��rIf�����?���3,6���9�CIlE��($���]���Gj6�"�$����2G*g�����Ka�?Lzd|)�����w�q"4����̩����-�.2=���2:6�4բ�}�I��(�t�N����8|��c�:��hl�Ŵ�#.D��%L1�[�ȋ���������~��s��U���ww=��qh>�#���ԏ%�⊤riw
�����/���MI�ew���z��c�^�|��g���{Jq�>�EU���该����%�$#;����fNZ�FJvN��Yj-*�B�H�����mOa���Ա=��O��#h�,��:*���#�!U���!�a�c��ڤ�`�ʌ(�1H��j{(韎<5o����������d�����J�ܦ�R��Ղ��%0�SW�[`�Y�Ӵ±��ܓ����������X���iի?��W�b.\�#����A/9�v���L�hu�꠳&���:��FS#�0aX� �9xr��������y=J�l�WN��w3z�p2o���K����ǰ���PwB�E����Bx�#Ms
�#�� &n��!Wk���}`��E��dJ��paݴ�
����+LZ�*y.��f�"r�]GƄ"d��r��YK᫼(��0��a��N�Յ�ss���[�ZHl�BP0�G���}K+z\A:>�0�G�8~x �T���e�%tx+��<��[�����^���	3':����E�*s'���8SAԄ#�y𲈦�w�D���!��G����ɕ���}��n�'� k�h�cEB㕡�Us6����G���$O� �R-|(�	�f�g�;!@�)㯼$�rPp���)�]���̤���g�|4ӫ����}���*���?��yɩ$�7�x�w���(r�����p�`G�o�d�������Iwd<)���ǘl�&=��yìTc�}*�uN�
��e$.�0`��9}��눧2���S꫹sW�0c�`��������������49��i� n~t�4U��	���[�|���?�A�q���Q�dz�M x�&���e�V5)q��pljݝ𳢡��'=��o��8��}�gḣL~�m���9C�ݥMBH2:�y�{=�	��K8���y麉�D�=�4TIP��=�m��o���N��E\��
+5O��j���M?� �2X�3�G=�S�^�Z�?���xtRfǦ���G��S���Hhx��;�����|� 8����E�b~}s{-�M��i��9aǵc��}-[>S!�?_|>�����0A1��홁IQTM�u�QXm;2����.ܼ�RO�W�!���	�I��R���7�'G�A���1��Н.krjV�����OK�*:?����	�`K1��Ç4�^�k����>}<�����7,z0g2��5;[�+=;+����ɝ \�Lv�g���c�gv�ޱ�|?���ĐF,�׭��P�.���c%�b������9�-�F$̀x�-�P��G���T�+?�P���Q��B$[����i#�dEN����q� �o�j|k����VD]��:�jh�n����������P�$x�F<%j�A�_�L���@�A������`\C��hp���E>O�LIX)�uppձf5=],�t8��ZC1<���^Q��c����V��:BJ�d��p{�)�K�-�l$E\$!6��5wUҏ�i���n�"6_3|<�hr����Hk�{i�S��=B���L!ըq��5Q9Y�a��Jmk	"������"���b�ݦrJ���>e߂�/j+��gK^� g�@�9&;�Z~.��PH���=)).ﯔ����U�=��9� \����=�hOǕ�����'*��q�M�Hlw��G�2`rD��q�8����	J�Ft���v>������������2��޾~��|�k���8lW�X}̌<��fw���
����!��$>j>��Wӝ*?�����9�Ga7�/��缁6��!��(~|6bXq܇^����!��(U�J�n��<h:���#~��'�̚�$k��I��OF���"�բZV�^:���h��]���y��n��P��~��ˬ7�=�/��G^�^���N����cʭ0�����m�i�0�WJ�s�����x�P3� ]Z�ۀ�;����s,�$��?0 ����rʻ��<�W�w�[��=L������P�U� �,���"�sW|�P�[�s6�V�@�>
z2��(e���� �J#߹���~���3��?Lk��o�l���׎��W�{�+��&-;�)��t��?b����ō�đem�w.D*g%~ǽ
.kYζ�	����Ը^o(쟍A>��i����`���������H��0�Xѻ�&/[���ԧT7ʰ��Ci!���/c�v�gV[%a����#��-�࣪ߚ�p�P%���+#�dE�m������ҍ��W�w?�`O��-�&P�z
�|A�n\ߖACߨ83�=6|ê�M&#���g`�����l��Q��!�r�V�a&E����VB�c�hm���rΟ��vs1�-s�����~Xd�K��Ƙ��2F�݀�����u�.>6�����#L���6֏�6O�\�u8{�փB+�7�]����?���Z�F�A�QݘF�4a�ۤ׾�x
Tz�=L:��������j�����33�/��z,^C>�'w7�/-��,����(���'���ms�T�n�:�v#T5'�xb���ǚx2�aw��GQҘH=n��+�;�
f��N�Z��Vm>�ȱ<ˏR9_�,�ώ���m��W��"�(�S���]���f��Q��/8�F[�N�J�vR�����wq�]U�����^9���s������K�sI3���x����h?��E%�4�JP֚�G﶐,r�z`��'��5%��Π#z�D���-\�����p��X�F0�%�;�&ňز�FMSo�}�~�� A8���$ӟ��V�e�"+$���7o���6W�����_�o����J��R��U#_���£��m��{y��f��*�XXF�x[5�8w�	%)��Z��'.dN�Gg�E��eu���|n�{��%���ǎk����{�Q�lB�j㷮Y�vͲ��e�׽|��ó�X����/�-��w���Fje�T����H���J����S+�[�;�E����wS/�O�5��5$�z��F{k�͒��*A3��)Յ���3J��,ײ�c̸�4 F�'��o�V���s8oV+؁���FlÖ��5�4�u	ڵ�O�qF�c����ro��^!T>���tR���P�G͘�OY���d��"�����R}�s	;Uc�l��Sdf�"�`���ʙ��U��"0D^���2i��ҶN�ѐî�5��e�:?8����-�[�X_��tW0c_��]����jQ�z�o�+�M��]9��±�U2���3U�_փ.{<O۰Ê�&��^v�]d��.)RB���[�i�z����
(c����R\�1�]c��f}{罘��4��9:;�Ze����\�i�ωA�M�u/mZm����r{��g��
���Y ���CF˙���H��M�ޕ���'��k?�'��IKԫ7��=L�`�+��KV��F$�u?�^"�[�e�>���W��{�yw9�Q�˘3)��эig��~t@{3+::tʎҁ�j��=u?�iw�ʾ����ݼ_��טH9q�K۫%���|�� �3������w����+�2?R���=�K��&����ح+^j�X����._9=�b-8X�������_��t��J��ثsQ�@�j�[���$ݭJ.D��=4�!�^W��u����?gf�;�zl�u��h�$�Wd��M*��z�?� �o�Þ�|E;>�}y�l��G�R��e'�u�M }��	4k��G7$:���"�h�"4��8�4{1�9�J���>������������=����V�_�:��v�"����rik�X;f���Ĵ�P$)GHu���5��2�%�|Ɍ;a��|N&#v]x�ŸLci	�-��jc��4��(��mQkt�eOd��u��`��J��7�_4�;l_g�;�b����Ou�?���V7"y�v�����.�t��ϊ�&�8����y$;$y��Y��h�:������D*-����s�-�8��W�=V��_����x�0�C�Ϣ�u��Qn��I��<S/�2P�A�����&�|X�K��hb�y�V���!������l�+�*Y�����%X9{y������5�X�Z�-�kuZ뤼�m�V�룻�_^�q#��>�.vf_�<)��ƚK.d��'�/e����knu�Y'�9PT��31ȓSU�{��\ C=^�b�z����İOl�ہ��2�<J�]�_�Om�����h�O" ��u)���9�UO%�g��^��f�֧�ܼ�_#	`A��E�I7e���Ͷn�oفirU"Ɠ`������H0�V��i�Q��'�,��c~�����=�S-ϸ/�u_ko��d7v+�(s{��
�w5×\��Rϥ��a+d��{�����}�YU��/3��Ņ���3d	���-qɮ����*��3N���s	9��ӄ�vY���uA�K`I��B|`���7�{�����|��hR(�f��qQ�"���}b?p1Ew��X��n��VZ������̛���#x ��]l�FN�	-�xn�w���Hݸ�ߪ���PA5"m�=�2<�և_�^Y�u~&��K�9�O�����=�F�@ �g�Q}~���l�5�����]G�O�͠�>�&��;�x�A..�֯���V��o�hH�e Η�k٬��?��9Q0�Z��?W�r�E�;}U�[�ܵ��F��r_�G֌���7ս����!m�X��C��� M
��ۯڝ6@c�\�k�؏���v���ە�>6����RN���7��5H&;���+#y-r`Qi8;~��P=�����qP]��}n(�M���o���L>�.��R�}���<�[R��T��m��ҖL�dP���mp�K��]�.�vU��WLb��b6#秹�߱.*6D��lƍP�0�ʕ��i��� ne���r�l�����J���y����nm��7jl�/��O����U�=�$lV�N�}�j����m�����[����&�[	ඞ�~Gw��DM����l��~L;�V���6�s1S��v	d_d43��Oo:<d��7����-�*�{QH���w�~���O�$����C��k��FD�r�݂��+��LY���,$>ckܷ�ګDe�1͑7J�R�rDdʪ*��㯓����5׮��|Д{Ҩ��W-�NjJ�&щ��WFF������,6��ug�x��1���F.P����m���Zn��Z����es'd	�$È�w@��PF�����m����9��*�����d�����W:r^���iۥ��+z[JӮk�h��Ӑ�ok��< ��1�@����$o��zF°y0�0ũ��C��p`�R"�4�'hN>���g>������z���ԋy�M=
`���#�����.�y�������$KIS�4TSOn�k_(1}��J��U,/�t���]joX�EcquK\E���]���%���	���.�#l�s�(�ͳ��W��hBh�SJCS�-t��i��B�g���nѽX�j~����WC?���5c3�e���bоv�B�#���$?W��Tto�{�uE�K�,��r
�~�P��Q�?��DT`�m�UVz C
�کW�`j�q�QJ��Cs7�I~%n��*!����.e�Nx���p42\���k����)��"���iF�{j~��=�2�;�.s����Fd��5�;-'��t[r��-ɯ]�w����'��"k�DY	��z'�n�n��S/�71��`�X�CV[Ս���,Ҽ️!i���N˧��V��|��lK�3���\tC$�Uv�q&ԛ���2G��?Ao���[�ߗ�{�Pl��O���E�^dv��G{��XX�R$}��LOn7��Fg#�h+!'c̷.3���_���d7����T�c�D���+�kP;��ҟV����^k2o]�^���)-ns} �?��/��8"q���Fó�M��ڼ�N�G�e���ȧ�-phJ~/���1���^v�f���mL�<%�@z�_�9���P�`3�)��Y�A��B`�n}Ê�6/YY��Z�L�D�M�c�G���5�J	�0;�]�1jw,̥�d��F\m����a���?�!	�6�k]�m7�7-?![����b�i��DK>��?1σ�����G�e���o(���&�<f��W�ϟ7��ߍjf2+�d�s�4�I7J+�moxhUP�o��	��#�}m.Ĕ�>f%�����Uu�%�T�h�_{$?L������=�.������b�n�Y�e���N'��,���٬Rǟ��0�9��_7^�*�)7�[p�eaAΟ%���K�rɐ��)�b�3 �}���#g���[�֥P����$�RPM��r�c&x��KU�ʥ���~��.�n֘C����`Ԍ$���q4w�G&{SO��7`XD��>X�68��e�S�<BWC3�Q�B놋�)��� �kD���iܶ���
�V�q<���+� ��������R��#U�1�%�c�9��-d��QywO&L�9e�xJf�G.��{g����+�Z�U��ׁG�̮�~�or�����9�ػ��0����=�f?�mH�<��R5�����w�6Hq>�F_�b�_HǼpD�9 ;�X)y�#iQ��2���F��X)#��=��	�.��;UT�Ei	����<�]�S7�ւ�*��2M��W�&�`n�TK{��8[��E/�~#2�9F���J(n�0?�u��5-����'�|o9������酧���s'��k�3�,���>0�g��3�.�o+��<��H���}��M���6>��1��/� ����C��j�O�Ed�l�����UK�uQ�n�������oR�gf�3��H��/HJ�y������;,��3Ԣ��;p	)[A=�CkBn�}��O\���\7��ƖS������m웶*�� �6����������܄�X��n1�Y�.u�߸ԥ)r��6��O�W�~�� *��k"��h"8(Z�wPr��JP+&(��(�d��'Xm�� Q�0�n/��D�����jcD���2WcM�r�z|@��w��io,xu�N��ҳ��NY�v� ?���g ���"�Z"Θ��]NZ5�����uܠY{�ў��[����;�O��St�4�s}��ܪ�G��:��:42�{��.�ݍX�?��g���^�\奈ˀ������3Y������zY���J=Ƿ||�떽�s<v"�
�� <�֤#~O��JT�/�����"6nV��UF�B��\�?j��[�Y\��UX�iЗ�	N�~�/������f��{�ڴ�5�����Ǵ��mOm�/({��8��%��x{��P�}��$��w���\�22�Z��X7��=GIM�G����hv���b?%�j�_}}G�i��j���ݥ�������kBq�r�:��oBF��R>IFشv�*rǛ�]BY,M����ؕ-�$F}�����`���(�\<�ܘG��G{qiY��{��Ve��|��۝g��n,��ys��8u�����F�S���͠���ihl^�(�t�H�MJn�t�ƶ~�/*0勫yuhd�b�ۥM��;4/����bg�_�V����nH�� ���7�¬�|�,'Ä�	/�RS6#�NS{��ot�ě^,i�?�g�&"�i�#����"u ������-�oc�dԻ{�3��������gN/\*s[.�NI�&�g�tgEDyL~]�x���� ���|��U�e,\�Y�p�eR���o���]7M"�:;Q	��ޝ�Ӡ�:{Ũ��� �횏�k�7ʴcm3��t��p�1��s���6\�| s�Cw���:.W�3�)f׊�N�y��f�p`��t�"�ؿ<�yku�L8�a/V
�(���o+��EVy�������\S%Z�+��B��h(�����|�&R�J����S����J[��Vtyk�c�#/C����R��򋊳�������f���H8|����09��i���~z\����刻Pi��V8����vT�����>�ZJ_<jf|2[����G���;�'�"-��Wq��Pq"ߜ���e2�K�>~��A��*�H��,��,�����[\/�y�Ѻ�����������R����8m�Yy�������#Ӵ���b*8��-|s}��A�~�?v�ց��-��Q����o�����L:kU��_v�\i<�<�b�:����1!�����~F�f�Zi��8ƕ�`�j+p��ۙ8�5���%�xd���}�z{{͏��F&�q'2rU8�ߏ�?�7xU�R��([�//��X�fV^Ah:䎪������9��w���c��^äѤ� ���~pPu�;��[���{=��/������!E�Ǖ�����E����,Rw95���DsU�B��B�3?n�H=��bd<*�UCI�����:+�=�4���2\Yu-�3q�m;a��	.�[I�������<�f�����2��3Sk�w���G�3�/ ��à}I�M�����x����)������K%��FdƭPII��$[L����Uv��e_B���(kSc_3��:�c��9}�m|=�z�9��~-����~�^'/jj�x0O��`�Y&��E�"'�m<�͊WK{[����ZY���Zr�eד�Ξ�f�)E#��s��Ӂ"�?|�w qp8�P�<m��<�/0�G����k����]ΊFؽZmPR�^�������	�+[�|��A�Vk2�ɜ���S�+ݢ��j;׭�d�Ю��'P��@�w|t�l�� �v� +b��_���	+���Ye��S_Y�eWz
*��$����_@r�1m܇p���/6rP�{��]Z�d0��:��J:eQ��s6��m�x8q�?��gf�b���g�ˡ�x�ϥ��O�B>(q��H3�DAIk��K����߽M�J��ge�7��Y�W;��f�@���>��*��k0�hefsvݏ@��CU>�6�>�5�g=��c�;T5����F�a��~N�ܫ�*�6��yx9g5�Wy�9n�6�R��\P��պi�ܿ�.D��J��m��hA2{Q@�Or29��`�Od��~�DE�ȗ��xxh(��DR0;o�E?�c�:]�V6�ｌT`a�����5��N���9j��_�nUߵ�9��yvBO%���ߗ����?�M��QDR�\���# ?�F�(�餒nj�C��c|3��ź]@�����H�o]o�V7��$W��P6ϵ��� a�f2��OG���ǹv��ח����'NK�˛�x�o����^�C4����[����>�gm���S����B�o��I���2�Q�ވw��3U�ϗ���
+��J�<ڭo1i���,��$"w-T�HU�������	���Xg�U�B �6������<��\�b �Y�=n�!���P9��Dg�V����.�5ȱ�����A���|c��~ab}^WH���yo�i�T�$-��gy#m����v�1^N���Ku���(q��y�좘���P���l���Dd}jj�[�ֺ�� ���J�x�b�d˫ ÏS�w���G
Գ,s��Nw�����dIξ����f�<:s��zk���t�J��d�;C`�t޷}���XU'	��m��Ʒ��T�O<	!���y��<kF�l���o�n�$� 'O�X��N�{��Ȑ�v��,����U��D_���&nњ�CZ��p۴��/�dP�`�����=}�q;�+�p䫠v��2zgm��+��0`Oi�ܓ��`�O|�GӒIZ<AE�&P[Y��;�]��/]��	L��4����okȘ~�
�!�d��ݿ�"-}h�6�D���"��I���%e/��5����/\_n=!@K��m^\�X+�s�6Y�GZZZ�Բ��3������{_������Z"�"gfvޟ����4P���w<21�J��v��=f�r��K��o,�Ϝ�{O��t3]x�������v��{ۯ��<�'i=Ruy�>s7xm��Y�R#ױ���4�J�y��$p�J�3;oD~��]�"5�Ɩ��A�([�bf�'S��N3Ή�cc�F�r�o��]Ui;A��Yk�Ϯ6D־�C���<$gо�����;��̕+�B޹�d.H"�d��n�w����,�f�o���O����c���@Q&�*"
{YFkQ�bo�s�b���'�W�3#�����oh�]��P���H�ߔ�<��{��B�"�Y�����r�nTW�y~�qr�4�#[�pg��mt1k�1iϕD���'���O ���HW��uWܧw����b:��<�9��JIߜ�k� ���H~fH|���}S%�Stg/�m�>Q�	�h^D�s�~�.���@�u��ՄOϷ�4}�5�R�~M\��dp>؛%Bt�T��<7�j��V	r,��J���
�uo�!Iμ
t��@��h�.\�3����!�����L��B\��$�f�4I�[x}��B�{�\� _���WEUV����g�-��:��jJd�qc�!��c�X+3���������)|�G����/[�ͷ��qp�nA����\+��NG)�����i竀����v�'��
��=K/TOܼY3e����'k����%��)�nR�G�+{U�ʯ��PyY�R^��(2�rX�Eۿ���'at�'�]X]�
���X�
:�\d�;���{)��1�D B�9Q;Y�߸2j׶���G�*��3p���&�3sm��睛WdMo�`�me�-'D�� *�\�;���������5r��1?��#�ٴ�v�����܌-��a1q���M��}O��m�����bWd��S�u{�G����B(��� zN�2��dĥ.�"���f:v����.�ο`������j��T��	(���Uầx�G^��<z��ޝғ�tKx�&/ѫ)E�����m�U;@Mf���m:�E�o0�������B �͕uw��b7�`*�F���W���6�N5?��P��#5�uKV��i�"`q��d���� Vq*`������JI �Qvk�$�>ڒ�%VN-���R�^�_��Y-�O���]ߢP���������+k��F1�`vkֽo/KK/W�Y����Z��[8]k��6{M�VbF|l��zJ���l� ������!Y� �fr�S�x,f�U:&T�Sעuv7�b���(gƩ���TOk��]�)�ڹvt���N�1���	�\8w��Kƍ����ȓ Oċ�=ri4rp��Q0t؏Ji'��ИǮ_��
6��'k ��*���u\&���0�Q�s��
gW�[�г�B�"өyHs�5�9:�3,��qXOMQt�faT~�6�j��[�:���W�E^yݣ�@no�`����J>^��>�pO����'8-W��=k��>��;~���D"��|���%Y���&�����Er���^b�}�T�d�e�~��V��J[zwu-�e���8���qxl�_9^@��-A@LK@��l*DUKZg��MI�|�`���$��x���Ċ1�H����|%���4WA�5���p0����"�⼳Ra�n��w�u�;��:�r���L�*�a�?V������k���~
�P~�G�gU��LG5�_m��b%>�\CS��`P4��gP��i/	������_,�Qt��){�i�1pM��>�9���v�ĉQ]�E�<���-="}��dM���w$F�Z�,3�s���J��8��'�zm�`�VxQ��ʫ	
,?���>�ih0b`���Q�9�!�p��!�'�u���Xu�;
��ά�ҋ��l���� 1B��~jgV�!ndn'�,p_�t��HC
w �җ��TF|.bjW��ʣ�_/.������-y�=Նp�c�� ��[<��̾����Оw�,u$���e 1��չL~[���b��o��"lVg�ܓB^��'�_�H{�{�+���`n��}ҍ�8���-}��-�&}��x�F=�\�7���gf�E�K�϶�5�@W*�^��睂Ʋ�����f�S;�l���< ���5� �{ t�-?tH�]כō�$h7�ե�R-pߜ�S'��_���o.o�=ڲNQ���S�����b���A,{U�`�$kOt�y�_F�l&�rs�kD�d���Q�(#\�� :�)���A:�(W��D:oY���ib��.b���M�����D;5�]��7"�����g�sȍ�\Cn���ݶ������+��.�S_�Q��m��s�R�vA�a�s��wJJ�}����e\��琝A������-�7ߐ. ���btv��Nu�)>�A�%��}�O���^�!�Z��D��`������?zԎ-L\�l�cv�Q~�qr��ę��^��H�()�� �|ud?`��7��Vy@9����r�H�8?��eVmY����RD��"���!�Y��*���A�d t�|�b������<�������Ǽ�"��d:���`~q�-����?u�fÒH��r��\��2�Ā{�4���p���Z�M���FT�����H��m�0ˬU�BڻE��C�y�+8�J�(ѳ��~�U=����C��ץUUvn�^O��s�'yU�c�����{n�w����� V���y�u���1�3���1	3R�܉r���f.�q��c�_/�W~���<�z�S�r���,p�%�����끿"Īx>�o�)z���~�(�r�86jo`���6�4@Zth`k%n��(H�d��,��B�)��M�9L��,@��F�Q��)�`����t��gZp` G�D9��kr���q���H��%�Ȇ)hƻ�$�){}��`�q�y��[�r���<N\j��3�#7���ж�!��W��x=I��s�DxJ�D8H|h~�,`���pIg?��ʛW({	����ʠ�)j��m�&B%w�<��D5�'q0}m��r?�Ζ]�I��\�O�I�K5��4D��2��:��ʍPHne;���c����d�ߙl�/�;"[y�]��^��L��f+��}q���_�/`��$y���=o&��xmh�/d�X�������G�N�9K�	�|;]C`9���Yb\��,�*Gʠw��9�B,�^��+������o�W�C��8@�=���(&Ӏ��4�[�祻̄M�'TC�h.u+�v1It��2���Qm渵�~������
�l@�N�䨍�����������l��.��嶝-$�(ՠ�E�뒡6R��>��g"a"gxL�:�"B��.�)�Y����/ݠ���ZO��E�:D��UH	��?�K_���C>�=b�W�CC��`�(1��>N�.F)y���	�aǱ���͙΄�\1�d\1<��?����,�gj^Wùf2<{v�n��s`�c�"�x%�`>� J�������!�s����;�T�&z'������?yu7�s���e ;���^P�
�	��k���>��x�V�j���# I����Ho��Q�/Sh��|sA�9F��PS����&)��O�J|����/��b�K�ڂgc}%7Ϯ�֎B;��j6JfY�o�m������4���0�d���r���.n����ܚ�RŮ�e���L���n���L�n����X�]��F^zi�>Mr�<�k���'��7�>au�Ǿ7��p' �D-��C�׼���qG��?⋞�����Z[�//k^�/5\O�7�����J��Ǉ=-�<&;*���g�]��F�H���;�n����'g(�!�G�e1��Q��/҆8H�M�.���շ��ZY���O�����iv�<�oK�� �}WZ��E��q�	@�����1��@OLH� �·�.�u����)�hB��E��Ѐ��x�#^��~J�4���n��ه���� ߮-���s���$��a�i=W,ds�����u��������t}��$z�(	�3�`�Z��g^�����7G�RJ>_��؛�|�58ٗ�%�$sY���A����"�	��-��[6lKy|XLL�<G�S�c�Z�O=&�Kx<�(���L+K�}b�j�h>D��|<��Re��Np!AmFlR|����z�.gW�,ul�2ɪ7[�B 9�X/���p�D�'��]�G)d;Hٸ������&l�� b��瀚+�����uU�]�T�ߪ��_�E���E���$U_�W�0�s�t���x�����+gj�n�o�˧G�������,�i��J��ܸ�%������i�h�~X�&�A|�����[��}��N���W~�̎$�.\ƙ�X%4[�p�/�e��7���}�O� ��]�d���C��2��%#-]��u���I3�����s��eŖEm/��(��t�i��q�N���0BUO����f2�+<Mz��IvI���< k��A쵈[_�|d�pugc�pu�o�0������z�ŻP�1Y�M�k��nص�L�z.G�ua�� �z	����:'�����J�n^V��g���S�.E*t�MX�'����f�;`z��;m�-�EFmH���g��)��Ë�q��ݥ�+�Y*Ȫ�/�@�˿i��
E�V�6ͻV�O��!#N�*�']��[$�l�2��t�ĳ�v`GY8�f�-m6 N�4���Ch��;�3�z�8>�p1P������t�-FC�h��H����fv'tF|���f$��[�0q�jY�u6%�k��G�!Y7v䶢:���T���i�\��H]�!����}
�m-��l^���xm
�����*�rK�¨ۇG�H������ڜy�5��ܘZ����&�X�lb��9�/9�/�T����~�^���Y�}gIm��̡κ�B�y���㟫���9B�bX�a���1=!g(oJ\ .Dy\0)�����_��u#�a ��ο�W�
Ű�y���9w�`mR�[vd�i7�������0�CK祦m}|O�Tl�p6rr�(�8�E�
I8�����1��~�TyYk64�/���=r}�躁+v�W�<��Ũ���N�g�m�3�Yz�Q�E���FO��6�	+�MH���Rh���g�pB�"Q�E���j��/�u��3����v=K�,95?��ɜ��Zㅨp�#O�d��bF0�/����i���%t�֛������_�x��[�'��_�ލ��Ŧ��&��"�?ȥx��N=���f����B�$��wׇ\���(�_��p�WD���OB���t�ǱO!��-�pN�ھp�L�a�pb�ۅK��W�ˬ��,G����\w�$��{���D2c�ĩ	�ΰ���@�W��_\ۛ�{���q� ��Y�a�I`T;��c�����U�)#�=5Bsz��,�����,M0U38F�3�Iv����4�_<n��ϔ��<mnk�g�����	�M|_�YG���U#hn��R�6׳	��^ÚN��WJ�����Z��s����N�QY�~vd�z�{���&3`=�o�6�4��	l��'��� ո�ee}@=yQrAT"ڭ��2�Yk�4ۧ���a�VO;#��F�\8�_A'C9�]�~��������0����Gz2uZ��.[�.��Ns���f�Ȋ�w�������Y/"���������숺���L�{ Gɏy2	�`�G'7S(�֕�q�|&X./y��M�s 7�+�_����&�Ѕ��U��-�M�h��9	j��x��bt�v8�b��ฌ��ɷT��5���W��ή�������q�x��#z8�͕�M��j|�woL��lEK7�i��͌���],�}�˕��[7�zݣP�ܘ�����o�������`��5%2�`Q�b��۹y(���Z8r���0�?ZG��\�j5����(���ICW�%@uV����7ä$���%���`� mX��mE]-��p�$�'���Ǳ�U��XO�O�v�N�z|�B9�QM�	߽�}���C1��}zY������ھ�ע��ֆ���#~�\O���&�ͧ�v��������:�T�7�>;3*�������G��e��Ps:Pf�aP�U�F���Pv����j��D�V�4���7[���t��35�"�.���W^TIU�+C�<(�5����F	����qw�1�ƲK��S�e��Ү	\��������_��M�O�G4J�����U�m�L� bi�v5�I'o���·��4�c xZ|�6�%]��o��ՃnND�g�zɖ�a��k�uh�������z��m����i����]D`��ۮ��X���F�`�r�NA�h9a����>$�jcq��ʺ|��GX9���c��t�#�� �>a�g��72^��/�JJ=ڃX`|]��6�:-!���W��r!��e쟹�`�����t���\S3�ВZ{�D�Ͳ�ő����_m�\B�~�p���N�7�:��U������cR���R���9�zf�̫fS�t�."�wZ�)��.�5oeG�7�E�=�E��^��=�X�C��q{#g�j�X}��@���R|�5T*ST����������?�;�0�E�����e��h�����7=��yq�����¾�wm]9�`֣�㯥��5�?�[�".���0��8(��RU������W���h_	@�,IUa����^k×�6#����~�N�{�.���)�g��_�7��V��a�7��|-m�v]��Mh�BK}w���.�������of�c �Z�aS{q=6^���$���h�@/�]����k�6>���pE�BQv��9��#��]Hӡ���jr}j�5BK���J{y���c���Q-��ɰY���:i0��%��hN���xaU�+����� �v�����H�� }c������H�ڵ�:b�h�֛���R�z��L6��Np�f��ADu3�������v�g�)��R��������;�(9��vO$2[����55�x�腞�h�,�:Ũ�d��_q%_F�Z/� ����i�xmd��2�Z��n�r6��fQ�����,v�kk>��_�ߝ9~��?���l�ו(@�K��W��w�s_H��3}��3g�ǩ�=x<Wڋ]�<�煟���O���#�5c&�H�Ywc��a�	n)Ξ�ݔ�=}Xw���ag� �j"��6���J�#�-m���:q'�ͯA{��u�M"�`c�;�Z�����M��;��Ѣ���~$o��<��2��ݑ,y�n���`sf:�eE�j�9�����7�nN؅\��ж���,W*+��6U.�ˬZ-;y����B�W�,Zh#��_��o�4pȈ�l�Iv\�U��k�7�1k�/%]���EW��T%!��F����d���]!S��{�f&$�Z]�쳡���~�D�_�leIp�%��Q��X-;Hz!\Ի��^+��ĺ��� l�W���yZ4��ғ�ɸ�;M����C���ıCq�T�!�{ߢ�����PZ�(��S��1)��w-X2w.�y�Xf�@vX2͹v�?��E��e���~�y����R@y�B�_���=-m�M~�R�.-͞/���Ҩ�v��l�=��C��M�
��F�~��w����2����ik�F�p�N�\����=]��ϯSvka�ó�x?$���s"���4�NՀ�x�o� �x�
B����ٙ��v~��Fw���w���Gݛ�t���v��6H���h�S�����Sxy�k��.���)n�ʬGo
P�w�g���F��=ևv���ɐ܌�?wz���?�w��<�������1N���@��,3l����>|q����Q�א*E�}>U��'��u5���Q�����,�Di���BZ�m��N��"��|�m���]��1�Sչ"�M̘iuϊ�/��b�t�{���WvN~(�1v�5�~�1:���1��a�߶�"�6�KD�[���_���7�����ᡡ�l?O˛P�Kxf�g�,���ͯh�֍�]9��ѵS=�ӷ���<?�>"�_/��}"w�gs������G	�1��e�y*�v3��2U�*M������(3Ё���:�k6�_A��qت�?{^j��k<�&����t��񣤜�2����m�+������w�?��b{����Ps���R��B/�E5�P�y�t��n���(|��.��X=d�/�h�y핊k��F�����[&����r����'�7�Ϣӹ\�{ݘ�:\������n��,Jaq'��+�=�����Eݱ��s%�� �P_�\���8O<�ѯ2�F��1��R��O���V���3K>�8�՟�2X��k:-�,V�?ϻ��;�B�@E�ٕ��	>И���7��v��tb�(?�.Ȃ?O�<z�q��Z�[�{��e��^3���Hmۓ����B�ɆQ!d��X�܎*����҂ұ��F.aV���ԁ�M���5I�UN�-����_��Ɠ{���J�����j�T�gس���+������2�4j�<*?�{0)�����U=x��}���(�A�Th~-[�ԣ#��fȟ�%G��e�f��$�5j���]z�����#7:S�ə����C�A��M--�̳+���|�&+���9�e���/9 4/�ʋ�2=u��<`�@	��#��{3bc�E��;�Ԫ�(��,�5�k�Z�b�"�
���$!?5�o�Ϡg��Θ{�_ĩf��`S�Wla��-��_سk_=$�+����H��3ׯ�N�!2��D��B#��2�l���J��n�����mD �dYsn�[����J��h?oC%�튥db��K�l���X��+e^��'���\��%�oÖ��ι�����(������h�Iff�H����qt����|]�z���]Y�F�B�Z�ttƬkzN�����T�DԐ�&�b�s��<΁�bj:���fn6��;�q�,�7-qa,@S�	� ���h���_�ܻ�'cgcZ�͔ ���$�CC����JՎ,����\��`s���+�E	�̠��S�_�<(��w��w�6�^e?x~�9oj����1��ӑ���n��{������e�tB.2 ^_��!sU)�}�诡���K&��7w���i�o<6�nC��,Ce}���h��SC,r�ˑ�u������t�c��ݸ�W7�����K�{]�V���̊��܆���1������o�(#�iNp�};���ݶm�/��2�ZMfPZ�I�(� z��hV� 5�t���ANs���~:Z��p�c�6��,�@0�%$��X �����b��C��8��G�-�ؓ N�	^0@)�`&��c�e`&}Q���w��5��B��{y�)��tb�������AbJ�/���
?���{����?(C[4sfh�����b�pQU� �}C=f�u0��N��7�"�غ:��Š_s��鶈��S,��Y��O0�=�A�mP!�^�?�V%l�0������emp�7��I��k�>NL�I-6���E��y�/�t3�G��ƅ�������<�нzJ�`�3��ه�������5ۥ�O�-�#U���-��]�uˡ�#�� W6H����(E����I_FA����A����_0���I�o�=�|d\q�������K8��������_i�'��v��T�k�3<�(�x�j��1c��GG+���h�+Ԇ_���<��4Td𱋵>;ռZ̋��xN!�Ty�ק�c#ț�\�� �Ƥ���3p�2��f�����u��T��.[����Λ�)xEi��ذ�h����%ʮ��ɮ�i�'53"��9�p����af>15s^��-�A!�^PL|��1�-�lr	m�?�P�Y�`�6~���:���Rg�\}i�v�u����Z/b���k��Eif.f�
��8�T�xrn.�fWU26���ܗps����`��= �U!����QQC�r�§"����ٺB>���;�QiJu�[QF�z��h���)�ß���,^�*%�O+�����) �O����J-��A��(���#M���,y�/�tz��*:|`�1���nXY �5X�J��Q�C��X�A�������j��V�K^��5�A)����n/��>�l'���`��>�q����"���A�0�-C|@#�� xmGkV���#3~��x�laD�0�k�'����g����߲�8�'�+�D�|�>�r ������#r��.r�����nگ!(���e�@AD����_-b�^�q�0�����9
%B�*J)�롟�7��	5��F����CT&��u@��4��R!�|��������^~@y�B������K���G+<�R�\̬W�w�3#��I��r�.y_r��8����� �G�����M�fI�|\(���o��٨[',E���_�#����BCQ���/��[�Iwܜp.%�}zIaf.�ȍ�:ڗ5�ZZ@S�O>�@�}��|as��s5����ql�H/<������c��A��JZ�5X>ػet�I��kC�|����p�2�����Ș:o������D}G�;�����w-G�>�&�n��`tϯx�5���H��A��h���z^�q�?tv)�ǩVڜ��"�d��=���10
9�s,W2��ed�����W]��������0w^�C���;V�К����ށ��� ���嗽�j��H]�v��Į��8������p7s�E�P��+�I��7��ADlY�C�q�t�f5tb{q��of����/�N���8���|����"%:3b��0^k��?n"��>S������8.ZU�Q�6��}�4���'_q�f;X�R_IrB���f�����}��C�c+)��<G)��e�Tcq �Y����D��G���l8_�vO�?"���;!�d�|J����-mt�4�/oH���z��J�O���e�fed��������\Ǳ��mVtO��Ռ�� �ة�.���ug�49t������*a������LS8�
CXI�\߳����K3_�z?�,^Y�z��b� Qɺ�ow�]W���"��*U B�	��=;��SYI7m�_�i1��(��SV�����ru�*��x��<��zܺH;wlZ��?b3$����F�HT�x��H��\|1=���9|�B�y����ʱ#���:2{蟻�
����dG��G\�ܛe|�ɡ���f�U����G�iM��ӿ,��7 ����Om2��)���-�΢��V]���Q��<��������|*�8�`P��=u��gm�z��y~�@M�ibV�ֲ�'�K�B�g��C�\��:�q;p�4Z�j�E|f��s���"�C��i a@�d�.�N�C�Av�b�׾n�6�0O�ovz>*��&z���q����јO�Sx~�2�'��x~5��ג.jj]�(�fl���r���'/�}��ە�)�9_���D1�X)�$bn�p�+w���~̓
5�}7�H��_�-o©N�Ȧ�+��T���Rɺ*M��[b� yz.��+�/�≳��3�pjQ�����-���;]yEt�i��PIH�&�<yvȢT1���SN�j�rd�ĴT��o=74�}O���p.OK-]�*����j�Ë�B#<��-�$uǇ�]=-�(Y��4͵0���������+a�����2��q���r� �w����-��I�Nf�
(�M`�E#q"��#z�6���v��l���f�GA=�MY}rGl�?�P3_��|�t|�V���@��A>��K����Ҟ1�7�f֩� xɻ�>�'{	|���r�Kv"���w�<m)�.��y6cZ����~�(��$B_�7n�Ud'�7D�}Q�����%\,����<��7@�\��%i��(�Jſ5��Uj(�7p�]�����.��Ԕ�����#�ݙ����|s��Ł������s~~�lJ�F�E�ܵ
�H���3�6��s����IƫaL�"�ʷ�;�qFQܾ����r�s��|����y�T_���ޅa$b�����-�B;<�&��H��o33��Y���T�w��k��f��F��(���Ͳ�����f�H�G^ה��ͤ��G�+l|q��!*���`/�����B�c�Y��#"8���\'+�ޠYWU0�r�G�� mF䉘"<r=1Q_&3H��9�:�Z���ޜB�΋8�+>n�R�A�*��fRJ��ݦ;I �.��{�}6��2 �+U�^,k��Q y|�S���v��j��ޗ���"bѶ� �������E�A�kW��Ma���R!c=8��ef�~8 K*V+c���PC5s���?�����P�ͮ�'YA ]9�k̐'Ԓ(�u�M�b�\��C�@�+���6�t���%�-�N���C���K�]�gQ���͠� �����_+];�+1��҉B�(�C	��R08�M�K�N�+fN��2��8ϴ2O26�'�{~��vu
=�"!`�`#�5�П_ۜ�CW�C��z�}�-V�W��J�����Kr/��|T�Y���{trC���*a��p�l�-N��\!��"�A~~0O�h�Hxh����-H��aQ"F�hz�fVŃ+�/��0�Hr����̜��Fl���0@{2�dvTͭ�؛��|��n�.	!��u���::*ԭ�\�-�u���|R�T��%��vf�K��F�!!G�o>���cu�]�ё|�4 ��������A^���LLG-�0EB��EJ�;J�١vzn��t��˭?�6����t��r �]xZ�[��Cc������U�ÎS1��Uy5<Z���kG���� ������&�}	V�v	˾C0�[3��}C��r�q@��v����������Z{C��;����h�9}d������p|LVoѯKUKf��F�4U�"�SSNN.��d�� ��./�,�-v,�w0�`l>e(��_�Z}8�x��r������M���3GS�_m���6i��r��İ�=�+-�YCF)L}��/~�qK�Jјk��6C���_�eЕo��^|$�,�l���+S-�m�]��$yFZ>���T�S�az��'�;�b>G��R;h�pI�n��(���
2I�gwBQN(���8
@��N=T��j�Z�!\D'uV�% �cf��z���wV������cm}>~�[["�.�.q�����'$�n�tZ�q���\}����Y�v�ߧ�V�-��e@�nO��V�W=*��������l2Q�0z�ӂω��2I5}�`�v~q-���A+<?�)2)�3�w�H���8���Ȟ*ފ~F$���9�J��S����\���I�6����(_�便��@�Uh��M���h�E
��G앪�ԧ�4���թ	�����~l������=�iC}9Ġo�f���1��c-����#��i��mf	Z��S�.�j>���;e�՗h�m?���~�8�L�u��_��9�+�R>�]����g�Ƿ����v�o�dKK;��HA��2@��T�٥^�����H���˛����	����? �Pj�U��uS����,1��­��/MF�����@D��]qT�>1������ m�v@.rG.$U$f��K�0>����2E�щ���H�"Ƶ	}#�h~�2��iaN(lƇ���h�P�X[�Y��m��cajWHL���9�Y�tѻ2�z�ȅSY�6n6o�]�W���R�Nb�5����{5�^~}���V+��7CΝs�F��?�-*4�5���aL�׭� �����+�<&g���<��D��,�Kk�6��m��&Mo�0�$�_=�}	i��ك�*�^$֌/�TKn2In�Z�ڔ�lBj������M�����Vp�WB�za�O�����L\����ӌ_u�	Y��-����K���F'�M��"��3a�I�|m��[���|)��6,�1�X/��EsZl�>� ��}�GM[$��s,\a�ŎVΛG�-HN���X�֓���ID��Q�ۙ~�k����R=;S2Ѷ;>i�ҹ��c�� ��-DZ�Ng=��?�P���e�j��d����5s�^I�;@�mц�wG�Er̐�G0�����^��� ���5��T>�g�:r>���D`��lP9�^�Q?�Ro>�Lp 5Zf*+�|Y��7̘*��(�K���|.}Թc���� i���q���̗֊	��tdI#{��}p�������5��S�Ð�m�~����Y424Z��S��F��}����F�	ӿ�N�����Bf���th攟�{�"���ʄoU6�yZ�TXo��)c#$8"Yv��ɮ�W��f*j�*�~��ҽ]��B�ų��z�p�t*����>�I�%0W�uMz	N�+l���)�ێ���%�Jf��wՇ�3��3S����f�����J�C����\_��}��A���	��+}꙰�wGG���y�@DO8�0fP_(����t��N2V�0M�o���ޏ&��^Į�d^��f����Sd�#�o-�r�}�͠�L�$���Yha�]767_&9�,����P�.%�?'��M�H��p\�~������
��Hp
���>��{:��-c�x��s���i�6��ceD��gK���m��-��d@Dx��~���^=r���|���;x��^���B�@o���`��<��?$�ݿ�=�����<���*P��+�a,H�1�y�HVGn"�O.����}.���9fѥ�V��V�:^}'�"�����.T}a���;�Xw�͊
�k�T�4`�"���=�H��w3Z���?ɖ��s����.i����?!ð<����a�)�v�w�XT�~�[��S�c�0_}<����UԀ��ߖ���0)�R��>��l�B/Ԫ���E�IDhx�3��*�0p~��N�H����B�%�#M���+�_ ��tFo�Щre9��|���;zu>؉� ���>�;i����Lz�0�xo�̴��c�{�e��� �V�tNWG�W۵:c��ݿI�m�Kڣ�����;Ւ㲃�$9��䳦u�ן�RJ*kj��V��;������Zw�i�.D����U.iuO�d����J_��գ��쓡���bB5�u�D���N��1 +"B���2/���W��N!�4����H�t�����w���n�9�:>��_/��(_�& 8U�ER���ɦ�<8�=&��yg��2�������J�I|J@<�0���و��;l�j!թq>�^���t/i�^�/�u�҄5q��LAL�������U[�9I�ʁ��J���S�K�^�Է�b6�*̺�d��@E�c�$�AyeL��Z��Ӝm(�!"ĭ�Nߥ+�cW!}ݝ�o����(���{�t���l�F�t*8�� ���k4}���9V����ϵ�5@+c6��>�>�6X|�1�Ǝ�l1��_���U��uJ�^�x�=T������z�v:#���X�;7���l��+[�`�b��R yC��G-�+��Z�GE-���-�0!*��� '�֐���dw���xKs<40��\�}ЉA����l<�{���xk����ǥgH�^�}���*@�-a*���ۑi6ֽ��U�2#�`�5�Y5U�r�޼�/8J�=���9�2��C�W"_�2ҽ)��0�3&�� I _rՂ��b���=\D~FD�yG+ �Ug�ӳ��ϪU���R��=�[)7�˂�4���6�Q�u��x�>+3�������D㿯����s�����>��ꧨSK, ���b#�Pu1��O�'�E$ OQ����/ڬ1�T)����
pn/~�#A���f�6H��%U?����b��_q�u/��vS �T5J�.�=Y��k�f�*��2�����5�Dm�0ł���ҋ" 	M���&�$����H�z	�;QA�zBK(� $�v<������r]\"lf�^k�}�kf�l��Z� 5~�ϟ�_��jf	ٶZY�l�MX�8W��Q�&G,X�/[޽��#����c��>��	)\�#��_Z��/���a�y��Z�q�,�;Ce@��^r F����/���~&�g S�<	��"�"P>����d�I�`ֿɿ��Ss���Yb�)�f2)| G����w �����f�"g�P�`�����Kܟ�@\*t�"��s���Y:I��k`ɏ�B�e��Ao�& C�S���~u���4>�7�� -���JH?��.��~�ŹsWEN�d�:������W��3��6��X���^4ͤh�BM��ޅF���N2X/��l|�w����2���W�����k2W�"\�s*����k@��{A!��T�(��� EΖ�п�m��\�=_�1�@�iǆ$�w�G��~�G��Y8�p:�-�����Xu�%�ĳ��ٵ�]�~\��2I�74��v�d�)C~,���`Qh�;�c����к���|J�i9��V�v��A'I*ͬ	
���Ӻ���Z��f���nX�ȯ��~R}��rs�dM��WadU����z1p��.��X=�t _���恊�4�b���7���}��u����Pd��N�Y�TIǂN���Ӈ#���_��S��~��P����'4�>�cB�J=:ס��:�10S�^�֐N�'�h�|��)w�5��7��:�F>�MJ�ro=��Ϟ<y��k���3�⧁sV���RR���7����]O�`,� st����ؘ���͚���!�+O�Q���!����:�	��ʽ�k�"��;�w8r~�2��TCKi������K�V{$i���Ai�Ղi��bCR�WF�*��g���y=�t�9ȏ[�5W�@%���g#3v�e��gX��JZ�:Noz�Qۺ;�GĦ�A�i17Q'�fZ{������x�UU~�B>=��E޿�1X	����#��kP^��n�6,bV%6�����&}Iw�:L3&���S��6�/�~[�yce��
��x���մ�Y@�:�t�$x[d����D���܏y�����-~ՓW;��R�uu�����O~>%P������������ApN��})��ݻ"��L��6Y��J�eŧׄ��}ȹiF66��F\ښ�A5�L
������e�n>�~��-zMwM_n���L�����^����L	��eӇ�N�;c���c�U�HM��zrM�-ԯ��<�l�	��`d.�f��I��x�+ N8(�ٻ�B���鉛��ɕ0chk-`��!�3�W�'i��%/린+�4��Y!@\F�##�;�����Ȼ�л����i�a3/IR���'
��U����<!���
�����ˇ���\�E?��B��Wj��],|Wf߯ƀ�Mr0�^Ȑ�g����<_�I����=����ho�G�!��8�}�a��I���6��dv�����6+��%n(m�i4��Q0��셁�'ų3p}�$�	�a�$M�O�-51�����֬�Ϭ�����;�����!�2$:K���I�D[�@�Ԙ��dg��#�6К��$2�|��F|H��Զ��3�c�IuSK�*Г����
r6�]�v�6MC��P�+E�ZZ�ڕ�U��X��2�?��	�W4ϟ�#���l�R��"���l$���2�\\I�%���~3�q~'�y^�&.K�li7����a?�e�μg�mt�T����}�8,�y3đ����N�`r�{�9Z�ܕX��ٚ��{�(]'�6��cc
��ހ�X���<���}逗�_PLR�$����Em�h�&$�_���_[���N�x�(���#��e����5��b��1�q��v�ɸ��0��d2��O2-lZ�ar���N��Ӱx�bͥ�;���лƮF�ղ<�ۮ�dڍ"s��pM�����8��nYz{<�����'��gG0��[g�ߑ�*M��T����	����2M�=2䭜�KWe�O�R,�-�B0)��޽�M^��c�����$O>`w&��N���#�fi~S�z�uɳ�6_@ 2Q�
��^z�NN�OI������ۆ69B������J�W�I�U7�M�t��sYħ��0�ZS�$�y���e4Wgz�${�P�d�F��p>mL��J�z<����v.�d�:M<<�Y���r���H<B�}M����|Ӭt�=�䫙 �s�`��dO2��H��qF���dA)����XS�~������[~��[���6]k�j�ى.��W���%w�zN�?�]���,x�a*N���`�:E+��g@��Hm�a�n�c�@m��Q#�BRGA�g��-�{��������*�my����� ����g�̢��3(Ȼ$V��-���oF�L\�vš��/%�ڵg�����X�����j���\ 6�Զ&w���n:��s���w{6R`D$�{�V1�$��OW�!��\�����(��Vۯbǵ��c2������*�	��':P���CYp|vwvV�e̜�\�ϖbX����o{p=�DRrj?mE�X���Lyj��g��MW��ց\������wƧل�C\�R!Z 	�P#����w�[E��|�<�L�R���w��η��p��id����$ucm��9���'��-F�# /����8 �j�Tϣm��'.������m'0=Z]��L��霛~Ҹ���VF�������i�fF���UXM9����H:E'�-|����z���;b��"�� ^>5� L���^���NZ�wfƵ�.$iwK��z C�;�V�]��z`L��)b�g����@iV�Z��[Z�*O�"�v��F���W��}c��~����-�au�X	�
��������5X[ۺY�-���(:�����E=��n�^�a�恞��%Ӹ�l04	��My)�x�:�7H8��z�ae�UG�Xƅ�ꪒ'xy�O���<��r��o�HN^�1Z�៮a�M$6,��7o�H9BXd,ܧH}Zz&�7w�����M�'�-��OÇ�:��q!H�n�=��8.�0�P�	u:d�����^Ư������l_���g�� �Y N��m�|����� @[��W���3ʉ'�v��@]V���3�n��ΪF������Hݼ)9�2>[��<K�F�F�òa3t~=$�輓���z-5�䗗Z�-�����{/�v��UN� ��555iȹ�(�d���Th�MB��or�j���ڶ*����5�Ş/�0J6f��&u7���vC̊CI��9Y�(SG�^%��v�D�j��М���[���ɚg�[��J#QA�7��<KQ�0K�:u%~K�a^�����z�2Z~.�ڈ��3��7���Lh6S��[�B:���Ś>�2\��dS�"Fuj m@@Io���W���n����{#g�=[|��,�g����[T��L�[�F�@�V������;=�/���t����z|���ӗ]��l�½.Q�S�΁�C�j@�_����A�	N-�εüeH����:-1�%�Q�:�Xo�r���lEv��v�hg�3�q�}�īÌW zƛ�7k�՝T��m�R�RYL�z@�QЯ���9|�@���#o8��B�`y�i���#�ѦN��2M>�x�iV����H�ٛ�/�g�s8Z��MS|�*� &����5�|�5�Վ���g��N��(.٦Z�ͪz��V�����H�t����K�k[؎1C�E�����E9�-�˽��7���;j�pn����i��W����݋U����*�$�}
aΠG���ⰛN�$o	�:��O��Z�VI4�!WHur�	
ىߨ�[�R�3�fa�Q�6j�f '�Zi?�b=8��MC�Y>ŏ��*c����+�UX^�`���ۙ���|�]�rq�phǩWu�_Oe�e�i�88��L�٢�Z1V�'F\�1�Ŝ�Y\�C<��Y�"��(w��h:<x�pH��g�a�����CE�
�;!�?�f���j�1N�B��*��!h��?�}�x�
M0�b�o6�e0��g��żU�h!�L�`C�(1{pAw��ڝW�+��赆�IS���(,�Կ6�f9�רb�C���cԛ#;3GE)A�����^\~K��S��	5�~ �b��`�d����,>wvTw� ��NXm��[ �[�Ҩ:G �7v4CNA��DWEYU\s�ũ���d�����=�y�p��_��(���q
kU��;��m%N:�s�� ���EG2<�1��f�&��a<��fc�\�C�?/����H?dP-���G�h��!ѝ�ҿ]���w�.���ș]2���J��	r��1��&S�Y�A�pis=G)��.~�Jd��.�g7�b�砕tw�[zx��斒�rt�&&���L9���G��X"�O@�N;�\gR 턉S�̿��c?����ޣgc���3�P�@���=7%�
ٟ���z p�-��*�(�s��~���N� v���+�rR�r��j�k��8���ɩ�2�u��o�~I�+3��/^����)�F�;� ������6�����Gm��ko$<bt�5�L�iw"+�w��^���
���a$D:��j����^͍D��HӑL"�d4E|�bD� /�rK��Ǐn%�[]WۅO�db�#w����oCe��Dy�ظ�W�W�+�q �fy�s�rw�$�L'�u�W�vZ�D=��;�?l�<X��=G�fa�t����{YC�.u�B�����W�.U���q%jY�)�p�jX�?�-�{�״�����4|zؑR�Y�9�]Pr�8|�{}~���u+;��J���g~L�M�P\h�'���{K��L�o�Z���������uV�}�;*�����G'傖���AWQG�Z��4g*�['EDo`o�<n��CT��,��ol�m�^ ��������s%[,���9��_�;���&eQ�^�G�����������`ڲi&��6�냮vTtQ��>X��)����Ւ���� &��w�TM��8zϚ�׳l�����A6y����+ul�{��\�1�c�a�ۮ�c(Y7	{�׽%`,i�p#1Rn����ڮ�+c����,s�DY�GA�8;��_�*%6�3�]ܰ��F�w�������ڼ[)���E><V#E�tB�e��~CY�YB���#� ��LmXS���[G#[�y����/�T��u���R�A�e�a���_i�e�|�O�����b�NH�x�U��*5	�����I��K�s��J%s���ʖrT�魰��=�1>zr�œ�#֞�h,�Z2�r�e>ߚkh3^�E~Q���RJ|�먚����L(�����\�Ip$���R�o<fC���!e݅���<���"W�&��Q!��7y� �s�}��B�U���w��X�;�e�Da��f\[���M�cPv��X�~�;�U��.�I�c\״��4����1F�JͿ��h&�/��}/jpگ^o�r�ۃ���T��*��u��3��kREfS����W�/m*\ўyPZ�A:����v��f��Y�B�LŋUb���~�+T���q���w�ŽU��ݏ"�[)V"�4��_Y$f�|���So��/�+�����1��ёX	���M�������U ����������F��pG����|�t�La�=��izqA�h�M���G����@֫��s�vXά��*���G�Mh��٣s@��Kݎ�_����-�.f�b8s�V�a��qW���V��O�s� �ܲ�w��j����wgj�O D�c����u�[�&�Z�G������{���u*��0%Fw��S"�}���+�����Į0?�9˞R�YF�Fz�*�栖5rR�`�-�Ȯ����}�p�R4�RN�gO�_Y�"�
�d� ��޸�����׿ U�>���C�.+�I7B�.�����]�}�ԧ�VZLqF6�1D�1?Y�]
n垐 �5�l�֭ �6�jU͑��쎌����|G�;R�IBs�Wl'tj�u�yc\���v��RQX��I+I5�M����4/v>tLix����D5��j٘6�_r>'n9W/5���z%)&����.<q�ߖ�����P["���X%��w�2mn��.��wZ��\�Oo3���n��m���4ur)���8���������Y�c�'�����+��A�O.�%\A��AR�/m>*�L�TE�	�<�q$T�lo����npk~Lϴ*/�@�o֮�c�S r9��+.�4W����gN��&\�#*��!�����ݧχ�ʐ��t��VK��ϯ 	Fb�&W>gʸ�u1-GC���G��f5�P�['�#}ؚ  �nyy0�+�b�O%ҕ<��
�{z���c��0��?6�>H-�Tp>W�;�B{V���Mޮр�@i�}��Z�+A�=Sm9u��D�Nm����$�H��}�k��t@�r��{�ؐ���>5��P�$�:t�W�o���v�/�����+$�zc�h�_�+q��.����,٫;?��� g�+������Ҋ�T
]�t��f4+(�g��r;��ɝ�C�*8ݛ���@�n���ǣ�I�"=ml(癭��qb�4�?ؖj���%�}��}/�ne�9�2��5=UOd������Pw,
2jF A�\�=���|� |���;=��͐�b���<@�]E��d㒑2!����9�u��0�M�B~�ƻ��в}��p4c�9��n�&<��1�U��z�P�H��p��.t��3�ePi�*�������iQ&�\����#��E�b%��Z h�<^������y���U�=)�
�0�6�%�2�[�CT#��B~���w���2eF�qw�������jV���-�V�>�_������+����I�n�������v��?� �2�q)f5&.	���96tq�*g�;;������)�Ml�4b�	�9f��[]%�%���ID~?�%��e��8O}��`�]Az�3�3=�4;��������䒉���>��w��ѥ��x���eU��W#xÌNgI�Qr�ԣ�Uݵ�S�T K��'`�rEV �ɩW��d�����ƣ���p��	�X�(�5�g��jJ��>�϶gӇ�L8ow�,?��%����T��o�h7�OX��M�/��忚2�)��b�&>�����7�?��rE�쾯Y�t��z��L��P�>�L�;�fZ���<����c�#&I G?Y�!R��^)�b��N_�2]�ͧ:��L���p��=�=!��
���8�$��RD�as�ײ�#52���6D�}%ί�F�YHw��e{�l6����n�<v��X��A�'/�; ����%Q-���Č]I;��Y��G^Wa��Df����6iY�o�eXJП�-�a6�Э�'+��:�OAߪ�߬q*�k+�ݶ�uoO��gw�<]a�l�����-�'�V��ma��/�&��l��S��D���J ܎$����m�޷�{o�I�n�4d���M	n�j�Q�a�У�!��B����߻j/=$�UC_z�R�fuA���؝px@�fm�NwQ䷻ש*��0s.!#lɰ=����������V���T�ظ[q(Uc5��m�A7z�}�4 ?�ͼb813�ԭs��9 �G�)�@��C��0�O��p��~'��y_�S�)�&a5t�=a�ʒ��][�S�[Z(C ���e��y� '<��n�WTn��ǌX�����1�B o*f��-� �X� _W����d]X��y��I��]�6�ڎ�	�JNį&�л~&����\�oԛ�伵q�}oߐ5y��,��)�S-�;8� 5�b�T�5����|��8*݅��u�m�@$���t�CZڳ��L,C�E�+�?��C�3��s�5J�	�J�`��S! �+���_��*�{t"�Fg,�FgB�����%MM0,�U�˂+L��OP\�r�9�5F��듷�֓;�������z�ɣ�@	�V3��i�x^A��[uQI�/��C_��]X����IL�C�=j�Һ�^t�&9��=���<݄�?ߘj]s4�6�7M�9b����[RPh���+�k��Ս�U� �Wz��6՘*T+6�a�}"�}��6��O���Mk{�'~��'�m�/t�^Q���'!A':��_�!w[%�A#r���Bfͭ��x5�e���'��G��k��]�+��QH���lmo�ֲ�<�~�}��>IL%,Ư\�v�&������}3�W< ✴=��͙����v�3�����!H�����⡜� Uv�<O� ��o����T��	q��V6����6O�Kh��HR�L��P˖�Ϛ9Q�����{�M���K}�2�~�-�ʑ,�}�c�N!��\q�6�((\����{�:t�%}9������DW'9͉L�4�є.��d�؞��U�l���l����n?[���\����> �]�7�LiF�0��7a����}0��A�p�I�tw��Ŝx�Z;���Ʈw%-�W�/��t�/��Z��F[�xG�.����KA��֜��I��w�W'=�ƫ�<�s����Kn�mS���P��֥d��R��B(f�bx�մ����ﺔ�J-�0Ei�R±ء��ė>��)KB�XT4
� �6[��,6u�_����gb���LY]%���U�h�p�U}��=5>9��~��k��Š�j�ְ;�������_&9�-Ƽ�om��x���o2Aeգk�%��F����%9��a�緹���·��<��|�6i��ء����g�+�UV�j�O�i)&���y�Cd�`����ne�7�e�:�M�Yeh�Oj�Y�*��������?�q���㶾�Z:I@Fvz�r]W�L�����i�m2���ք�~�^�i�o��)u��,5Uw,N>�HՖQ�8�C��Hl��a�L�����pT��U�`�$��h7Դ�܍�14h��-�@�B(E�Gy�#יD�{�$3��W�}�����o���R��=)Y�l�=R,Ax=�����#
m����o���	{�W�5'�2x�c_q��O�bx��F��u��9wy��-��c�A
?G1T���=7 �~�A���e���_���$�f��L�2��]����f���j�-�&[�X�}>`+�Ԑiz[q�f�a�p���{�����RM�)�W���l@��|wP4ZC�=2B�!g��Z\<��gDV��=,��'~��K�]���m�n����/ƽ��*
���M���7�������
���n���`7���'�^���Јa�4�ı�+�2�ٓ��G��`��U	����@�9�n���-#ҍb_����x���{H p7�_n1���������f���G���m*4<37u̼;�f�t�jBv���=�p�<l�Wm{��K�u�z��1�|���y�<�a��h�k�t.���Cbs� /��Ԑ�͍��� _[�-*�!�ӧ<x6��q�Z<�R�������r��X�ʹzvC�QW�d�C4laYs�Riy�i^��:Gn�:�o�͕I����?�0Q%פ�x�B��ۢ��H���7�Ÿc�zXrSا�2t����A�ɢgn&����:{�,�m�+���U]���B>Wqi�����q�jNE)�ڈȩ���
4�I#��ٖ7(+�ي�>.!lf�kQuߘ�����L�6S�.���Il\W@ij}[ ��%� �<?���-��&�q�oɷ_�~�0���f-x�ں��;>jc�\�X���x�vMǽ	Xtk+��0���t�.#���?"�J�{�R��D_A�x����f��n��5��5�=%@�'�!6`�0#[ ����%�����g�#S��4���(+�S�G�85����G�{��Ù=���ܠ�09�Q��<D�n�=��0ټA�|R�_x��-��,�NSC���e3S���U.�R��!%���/�6V����L�з/��Qm��#_t��u����TM�<�8�
���Q���=<�̝Ҧ��@D���3$��voəa�\�ٺ�����ʙ����`"l 聛���e��S7�* Db������*��azn���h������p�iL��'���Bۓݐv�g�5�^�>�W�F�,3㻠�:�!���$F�xL�&v�	 vZ^0 �U��.�ʁ�"�wp���}�Ԙz!�H;G%��4���Ia��ڍm��[��K���-�w+�P���v����6G솢�H�}#�=����@!�V���)��L�?��ۧ������%RyCi��l�9f�Ӻ��)��pg����J�Cxd>�ܗU�����(���CX��JRGϧps��"��~�7�5ɻq��{�|�)�B�c+-�MP���z�a
l��/A}�V�{8k#��
Ȓb���k�jn�Z������p�k�Ej%=���nPB��-����S�,�\]��Cc)m/<��,j�m�?�{z.�� ¬\�6���D0k�f6�#6�~��}6Rg-,犗7����-�{-;ɏ��-(l4��p�t o���}(I*4�,�4\���]��Q�a��HXn��V��
��~�g(H���E�U�b6�\�_�6i��-�e�`���)/msw��Mڔ���&݄t�W�����l�� +���)�
Ц!��Y[���S�U���_�r"�����b�|#/U�ׁ5����5>z�ю��4}��k����[���y��v��LC����k1V���[-�@�1ٛ����t����gm~dm�n��Š�aT��E?�j����������C��3���� �k�ʲ֭$�Jz�W���.���Ϳ�`<c�X��|&��|�G3�*R��7�6y{�?P�2_z6uu.M�j��u�n��fB����t���v��;\�17؟f^�Ì�~u�����3���7�J��m��w�����ZS���0��Ǧ�lK����R_
���"��y�Ց�:$���c�p���琇㐰 �K@0���-)^e�N�׋��%��Y|�a�K..I�P3�rK��.�a��V�S	)gЪ�ɓ��4�3��Bu�[�h�vl��i))��T��!�
��eXO�z��ND��Q��k��`�5��{`�l	L��w�B���\l���5y�v!w�e$Ow�Q<v3���hˢA2ܫ#n��\�2��N��l�{�'������w�I�/�0�P��a[�̋Y��.x�Ůi"e
?;�}�ȓ?���\Cr�r��i[�R����e�p��=�:e@��;�F�B�Z�8m�,sI�QG�b����}��*�p�W���I���Є��B�6�'���a����'o���d>������(<���FC]�㥥]{۔<$��K*�v�Y$���'�3"�e����X�#x,_~T�f8���eGGF
�K��;<��&��J4�&�J�Q�? ��?����=�̻)��]k�^�$�O�4���y�b������;jP��a�%��� ��y�>ީܒ�%%V<��p��<�xx!�,�@6I��>�Tǆz��&�������:���&��j���>���8���n��~�������+�<f/����-�����æ���x���G����pEUE���#�9 ]]>6��ld�"u��0��H�J�B��H]�᩺cA�����,y�M�	B�Y�A���RA�n�q4�`i��,�C�����n�tlM�&�`��rgT�8��y��i�ت�H���kl���Sf��Q {.h_ʝ���[C47Y��J����X���$�Z{q��ᚽߘ�<wgY��z3�(o%!�����������m��z~�t�)�@:��e����p�C��K�:�3��H�����e�umg��t�2�o�|������`�v�B�3z����]d��i����+����JuZ�	�A��4����&8���/��@U�{��D���Rx\k���*����-�<%�������j�,+�<���({s�j��k�ιm�6�ć;�5��X`�����B9�)�ŝ��2����7b��c��D�N��=]��#z�9Vs��cҦ2bq�q���ό�B��
�ޞ "n����:�h�^�8��-���;��
��Բ�~�HW�6����Dj�9'�&�YW�.��U�Ȥ�!�I�'��C�8	Ɛ�ކo{b�5h�Ì}�jB�,~�%$k�C����B� I�ձ�vH\�5'�e�W3�G�K�g�����~�>(�������L~w��aI�v��6�t�n�CB��-%��)K!�Z3	^��i����%�� ��-�QK�8i�;��1=oō��M"�{��g_&L���-c	�KF����U[!А{���կU5k��?}Gך�Ҕ䁒pf�ھg�8�i�����W�j�f�s�[���Сx((3	Gj�g�e�=5&�X��n���.��0�2�ߖj�47/C6�:��
�@5^���۬]�
�vҟ�۟��~Jb GB�S�g�|83ks����
Z+�����0Zn���u&ѥΫ΃|#B���w���t�k�����D��.���^�������s�[?@�^g�~�9ݩ��̨VE"�m�
5<=��`�h(�@t������g:MAq}��tf��n/�=��Н�YB��*=!� T�<�;�.�0��#!'��!����n�,�D������&���jȠ£'�4�i�IK-����zD��dmH�2F������>�c�ı=M�y�	�76�-�a����њ.������y��^�*7N�a�T�f�߫|�*�IC�"��Ul���7c՝ԦS��E#���Ke�
K.���]r�pK0{)G],�ŝq�!���G��~�ք7]k0 �P�ʗh����-��)b`0v�G�MY��}�,��>A,@��� �1	��8+��w���V�U���Et�5���/TkK`%X�"��]��hh՝�z,�1fX�����O.��H�ӓ-��;�G�t��f�o�t��e/¤8����r�Ҭ�.����UrS��4WwS��|��[&ێ�0��u:��yNH�釺�&���OW�5	\�������=��/�^�^0>�v��2�PHx�7��o[ո��ppY��╅��_U�������GE)�͌�\n�t�D(�1	fצ	o��RL���ә���1��o���C񉆟�l����GR�E��Pc��Q�Ҿ���dйt�0���C��>(�������b�DxxTt�*���}��n=�]49�Z-hnDޯ��c4[�k| �:��HRݝ�$E���6L��M3��m��m��X2�t�J|�j�z��'��*�n|����IL;D��_���0[��0z)�,�9鎈|
�G���x:�3X��Q�a�B���1����~�-��m���1�'��y�{$� d���uT-��f�g4*�='C>�ͺ5sI+��l�Сǌ�z#��}��rl7��"�l/o��|�� ���tK6���};�2@[�y��'�>Pz�1��z�|Z��OkZ9�!w-�@�t�N�R�/U������z`�Z�����l@d�
���#R�����C7 �t����G�����w�W�uɠ/|��e��7�Vrn��!*v�+���r�G��N�9

�#%7���F:�g$ 1�J��J]!IR��灋n��l��v��4�R��)��J�m��r������U�e����6S�9�((�]8+�q������� �eJ�@^��I�����ŠD�f�#�KB��I�p=�;����U�P�<�&`T�V д���.e��yv�����k��� ~���;��i����uSɵΘ7?O��*�JY���qQQ*���B,��z���6Ľ��\۱-"~I�,��������ݽ6�/�0t�Г?�2�gm������Π4��4��ߜ|�;�ݬ�����H�m�^ mz�1V��p�#�V�f��6�τI��:Qjb�5x�����2T�I)Jd�qɐ|�zw�\���"�R$�V��hK�8!w+N�(��]��U�����P�K�s��X
�1Ρ����w�?�}ˣ/���.�zrI��d�U@�O��{k��6*D�ͪ5�պ�B���qtpD��l�@��{�6�z���T��ya? Iy7���>���ϊ�3���l��r�Nbz+�	4éT6��L���RP�
O����Ҭ��
i�"C{���(6���Ŝ
J����єCJ�k�nq��޹i�.�p�B��:�J'�P�w�>���+�ses��˂M��?�T���u�^_Y}WOP\>q��'�H���iA��ܨ�&����o.S�?<�@�+�Ҳ��ɀ���h�m5)���SG4��[���B�o�;Q��p�.�i�!;�KԱ8~��_^I�g�������_<Hv�� � ���f�?��|hBh̜EiFY|c�;����)�J	 �������U�.U��J+hUM�햙^^F���Y�7ިa�4&�$JS��p�-�УUOP<{��hP�Z��1��s�#ot���"�͕��AT o\=��]�ס븏�l@����0��^�O�)��"���A=�5�E|t\�\�J��V�w ����x�Q��:�Fe(��Ĕ�������w�~�;6)"84D�����fV~�r�Vde0iZ� �)�u���[Ɖ� =�')>zJ>'����4a��ߌ��ޙ��v�Xd~D|��Y���R���Bb�3���W������6�*hS�U� �R��s�W�Ѫ9��31Y��!��R��8��`]��kh�A�����p��0�%{�mh9���w��~��C�yRNP�!�*:��xl�x�Rq��'�V���ct�®~������FAX��R3">�tg~J�4jR:X��dC�;#�q�Q7�ˏd��7�~�6�c��=�6r��dK�ٻ&�_�����J�o]/��Y*��F�;��}P.�dq��XТr��m�F���l�Ú˒=!i��@�[~bN�-HA���]b���턬b�s�:�"!H<5��ϝ�����:HuU�w�mz�V�S�YնS7�m���8`��X��:[t�Y���$��ܾ��X:w^y���ȝ����ڈ��M��3�R��e��r��8�r�P���(�|����V(��)�>�j�յ3qO(KG��9�=`9U���n���&��rJ�R�]|b6�(���3�]�q��ԫ�J����l@S"����Z4A�Ŗ��}:C!{����Vn�z�C�ug`N�)F3�_K�Y�k�R�G��L�U<JQi�z�,�n!zB�O_l��H�eht�;yCy�ƟH��^o]���p[v�vn��%�cƳ�7pE�_E�C��SuL���_�Z4�=�y��Y|2���Ƚ{�9K���_�u�9��+�t�+���	��~g��'Vȭ��c���\F� ��֔D���f`�1d�,��r~�$	Q$��ц8���{�A��vq��uW�J^�Ec����7�e4�
۱��T"���ʧ�xm����-m*5r�(X���ǯ�=�	�N���~�U|����9���>}��R�d��R33J�u��]��W�YI�G�vd3$+�*o�S���|J�\K���cv�:�:5(�Z׿��]0�l��,�<湥�Ņ�P�G����<J�� Z>W�rK�d��1�7����!*g@������Cƻ�3t�F�G���o�;թ �I@�یh�'�)��_)"�U|
,��H����[*���X5��>��9q
�8hR[;���tF"{�;6���p��������qW���Ñ�'�Z�b"�dz'�ߣ��R�zJ�n��Z��2]�8+p�-�ǻw���ƌ��a~��~���ҍƲzV1V�n~J��9�	��yz��{��Z�cM0>|X{����6��ϯx�W�8Aj�{2Ua���S���Pb�y�@W��/�a�Q�p#n`�p.��te����vtvN(���9���;�U���΃ס���)��xZ�8y<aC��r����lm�b��s'������6O�&�;�V2�2�K����|~�z6��>R�gV�%vb Gq�����0�={�Ǖ"S���SYU]!,ˉy��� c���u�=u�e�R3x=�zu�I,,���xhM�gT ��QT��z��g��m �:wܛj�m>ٛw)W�� Y^���9�o@�cV*.��D�|�M�A	���2ԁ�ɺ{��W��Mlc�To�Wa��g�$�.�;����<�I����dke���|Lull�?J��i�s��h>�w�'#�c��8��V���m���g���8�����Z^M��Y��PK   �u�X+���q6 X6 /   images/1f8ef630-8a1b-4a9b-bd39-2911f79a26d3.png %@ڿ�PNG

   IHDR   �     ;��   	pHYs  �  ��+  ��IDATx�ܽg��y%�V�0ӓ#�03�9G"�@0��H��$˔-��k{���w���?���l�eK�%J�$R�A 	"gr��{R箪{�[�@K���������;�y���O�7�l���a����7?�_��sw��{>�@<�խ�ہ ��p6���+l�^�&�����Ŀc9���/�X"�˛v$5��d��P��O%_�8��y�\ʓg<#��Ǘ�y\���g�~_��f��?q���f�o����x-���i���6_�����g�i#���P޾���l ڛ�9�I���o�+�����y���&M�e�*sV�/�?k'}����<>��~�2J=V$��c��_�t���X?~m����}�_��?��W�\>�Ϛ��۝���v>?n�y+kZ��Ӱ�i��l>m
~Xy���vд�e��6,ôMò�1���sY/�aZf7�,�lar1ø��o��/!�#^3k���@�>�-����%`�,�^��/b�^nq�^���}kv~���x�=��\��0�o����z'��4����kp�נ]0z-^��	1�v�m�6���MKl�����m�e������ß�8�ao���o�~x0n��all_�W���[��h��c<�搊�ҁ��
`4���8K�L�_fZ��	Y+�%��c0�/"A_q6`f^�֏_�Ɵ��S����Z���{B�����5K$$�Ɉ����[sYSr����_0�6L��_5��P�brJ8B�Ia��#��/"RgP=zg
q�t&�cL���q��~�8�q��Ka��$q���@{'���:��u�x�x����}��������^W�s�c��/���<����^���o�Ɲ6ۊ,�����+���z���{��v �oS���C�>����m���xG���w��A��'� ��ȋǏ~yL�y�@�	���c��$��X�;����q�`�z. ���'�U�|4d���k�~����X0
茟Kt��;k� &��g�<:��ὸ�N��1�},�ݲ�: *n��w 29,�L�˟|׷I r�k�Kl�~P�7���]�����31����	sǲvϳA&�6�kM�!��/�����9���s��`K�
�w�H'���u�|������3���x|���(��t���[ ��q�P[�5ms.�氎W[�8���lF�ě��o\珠�̽�����>	?� k���C7��O��P�xN�1�����4��np��׉�Il,:i�D^�^�	��Ce�(a��������̉3���@0�+˴]��r���e����Jvo��g؆c[���G����L���j-p��p�-�!�A�
�9&
����sMG�Y.�3��/����+S�uq��g�.0
�2��\`y��Y��ĵ�e��;ƞ��Sq�B����2i}]q ��9,�L>��Þ1���d�4�bJ(���1	��3קF�~��ί���~�ޡ�X��ӹ�b|��$֒��*[�an,+���5������|�>e�a����!s�u�郱j>��^0k(]��,~s`2�L�La�<�fXg�r_�
L � �l��Vv�+��O�f�L��6��`�˝�뤃�!�W�^�FM-�a8�(0(X�����������{�), ��m"�B��g�
Sh��_�P,�U!���23���������g>�+��1��^�̀�rxsI|�rP1v m|"�l;^*R���o�w���0�9P@ҙ����<����֋�,3@e%�I��s�X���Hڇ+���@��1�d
�px�cLL�#l݉3���s� �2 �`�3�wM�#��� �0Q�/?X� *�d9�0M��N{T��Ú�p�m��l�WY�n�!��qAm�� �ۼ�J5�c���'Gr�>��e(}����Yd\�j⬻4&������L��t�B�����~�a�r�,�-�q��<�2���X'Z(S�^�W���],|�E%��D`I�7=Y�be��E?�����lO��~�3�R?n���}M�&=�/��Ob�(DGVPg&�F��X��@
)�<6���<�:=�C��p28����*|++�y�0�l���7l�����/Ra̿{
�c�,���L��N��añ��-�����G���s�wm����2�	����cb�*��^�=2���*��r l��FAp\���X�Z|X����..���xd�4�R�8���D��%D��$�6e,�y��l��1��,㜙:y�M@=Ͻ+uX�h���l�o�y�@  ��tÛ)5<�z.`��4@��8��LB�iNhMy����H�HB�bP�Oz{{��@�����#���~o��8ޗ��T�I�\?�סy��թ�e��S r��w��x'D�C��A�G��
㻽2��^��ݯ�iuȣ�{��I�x� C��<.-�0�d(ל�Xw4��o������Ͱ���_u$
H���8Pl����8GN�|X�E�����o4�'�U�h�|��8E��hT��-�DJ�����r��%���/%���O�pp�p1��U� G�dC�V1��1M:�"�^z��.��L����O�^�0p�RɄ��J�~�S��a�òl�"4x�Lkl�*4>4)�����n9|�>vVn�uHI�$	G�e41j��:̢���$ԃt�p�Ga���T���c��P�X��i��Jo�n�m�&���Ý�� ����;BڍI����S�8w�P&<>")����A
ޘm��OjWA�y~����s�>��@�	�$�BK3
�E�M��u+��ˬ�i9�M�!�Xâ�f��5ˤ����<wQv��H���?j)��W�'�>p��i��׺7 [ V�9�JauNQ�g��%h��<�j�s+)���N�=>"���g�|L.�+��5226&cc#��������bQ�<��9v�|�_^��/K<9*�X4X@'�"؂fӀe��� ��ftյC�萉x�eO�t�x�n��+�vV�N�ug����,
�� ��|Ѽk������G���=a;_pP�ym���a��Zjw�ǹ�D@w=�R!k�S����h�3���ӓ��<��'�G�B��dhpP::aa�RRR"�ٴ�j��/E�e�fQ��Z�$����r�s@z�ú�3p��T�ɓ���G����qT�ՠ�^Ú����1�����\�l�<��2��I�����
�HQ��T*!�!�\���:Y�|�4Mk�����~����cyX�bu�rt��ry�k2�
�� [&\s��\3aV\3h��O����iw�s"Xy����a]w ｗ!�] �]^�]�|b[�,$�Ft>����Ї �����~�,	˗��)Ol�ո\�ňF��5� �:�J 
��2$1,�4��Jyt�RT�7�= ���$ϟ�����q�4�p���"��)m�kɩ��E} MR��Q�%��x�y��g���T��:%>0��r >��� �<yh&��IՒ��x��	ih�-�������%��I
,@���J�n����ʻ�8����tuK���,g�3�rw�~bB �S��Lù��~�w�nS���}�]Q'�j����x��ѯމ?�jA'Bܤ����d@M �m�Y0�o��1��t���R�>����Ѓ�����II������`<S��r���X���%`�ἍI��ɲd0<��ޡq�|3΀��Q�ɧ�{������ը9^�[�0����-R�TD��2��ACc�mttt���Y��f!��+���O6�[bl\=���))���6�ŋ���1�%	9.�Gׄz��8�E]k���"=n|���TUMx���a�����ٮ�n;����uK�g�s��*L��s���bH�t�6q��@ES,Ƅ�r��7�b�{���;�߲��pq�C3��\s��@�g���;�����v ȆS��~h\S�W�vt2M�9�L^�ǎ��R?u��_��Z�󐌍d@��c�-����Hag�lv��PçJ�'tYq)*��2c�f�Y�h��t��i ��p_�~��y��z�n��觐Ws�322���e����h�L9s��JQY���>\���.�bl�r�\���R!�li�ˍ�[n���L��d�B��`RL��u�?���Kw�։�;��r���Gv2��V�t��"�pڮZ�Yໜ���<&�eL}͞0;Ca0�,#>��r���M��JmeXn]����@GFF4��������h�<~� P���SK�Hb|P�++d��yr��5�W�D��N����	`��y]ٖ�&V�:��b? /5�e��<�aRrh������ ��9%� `�����ޠziIRm�V��?�%--�pa�T�J�C���bx�q3q�N��3����:u�0���x�0�8Ὃ|���q������g"
`��,h7$��4<�6��۪x���>������+$�E��]�����Y��=�b�� ��࿃tzrt�M)
zd���26��II�e||\���!"��I�L�9���jC�)`J��Q8i�2�hQ�4L�����r��[���a\C_O���X�rԐH�>�t"�~�_�`�PqHB>KfL�*��K_<��zn�A&��)��O���(�������1M�?q�Kk"�kgevK#�Z,}�qtdDJ�K�2��p�<N�	 {���u���lMk@� ��hJI���g����>���l&syGK2HI�Ĳ[���y�  V�N���aH���&�\�u�1��k5.G������^�S͐�[jڹ�l7 �Xs}l�D~���1��?�+؝$��;,ٔ%��c�S���0�V�cQJZ����B�%��F{�'wi1%g��g( ��^��W���|)\G�Ú#f]�'g[�#@n��37��4�L$c��46��%��y,���h��!x�����(�x�?��<4c.d�(&�<V���w���|V&�u��6��^𶕟ȩ�x/Nt,����7rM�臷�q���]ƪ��^MS�F3�Ҵ��=0����d����LjE�_'�r���\5��A����(͞ǫ�U��M�G� ��\�C��"�'��CeKM�ݓnrbf^W[:9U��
�Y5�x�7`h4�k|L����}z���@(�Xl��0ːf��9f�e{�5�^��f��B0���1�D�`>KS{�3����,{��9L\�1,�յ*�ѠhYT������TB�l�kD��9z[9]A���$�����c�[@ɄD5N�eJ(�o?z�qJ`
�C�Ƅ<n���j0�|'�U�L�Oi��,�g�B��"��T�'�Nb�3j�`�`�Q/�׏�Dc�RQV7����9NR��!u}F0I"�PD��1a]}}�70$�|J�K�2ɐI��%gsXpL�c,Bѐ$���@�cJI��:-� �_H��Zs"��QMib�X4�(�ǆ�!�-��Ӵ�i-;b�2s:NSk��aD�C��(�{�S-�����7	'��;y`��1o
��ܶ��ț�LF#��|�҉26�+-�Ϻ��	9�V�}0^mx^����|��3����f�懥-7mS(+�N�b6޴�����d�Qt΂Xu꣌,A���[�b�0iQ)LCEm���TȔI�RUQ	/) %�Q	��������:�_�Hč~{5?f�mwD'+���gs����Bc�S5�RRZ��x�� ���&���[z���`L"�R�W�o_�E��;�z�N�����yY7��,pq4��o`P�ɴ����<L[@�,]�Q3��4���h8ð�S�m���� )c,�C���%:p����p�}��{����<��M�xԃ�̤s��b��h�	�~'�a��a�M�[Ӝ��;	D&�S�NT<>"�� �ϧ�@K=lө�q,��D75'��+�AQx�o�ᠮ�DjTL�b�c*�&�E�jz�̘6Y&�U˴)uRp}^e�p0���&,RV�M͢�ӈ��(l,* ��*��3�K����J�2��$ ��GF�Z��'��c�r~���ё�1���;���.M��S`~����'��L�BR� e��C�ϰ�m�a� ��!���8���`��5eN���!�L���Qs4��u/�Z�OE�ᄞ��iik���YR	i���i�>�Xt��p0�,�uB]�����q�kNCd�~�Qyq����>��Ib��O!L�u��`�p�HM�͛7���&�R��x]>}��\��,��n�Q^�jZ��j��Wى�8��q���5����u�R
А�6JIq�����ҙ����.xA���xb����S��
�� D0'����⽪*+erm��~��Ur!��=����"��14����b��y`�Or��u9�zU��u��I���3�W/�-�qL�3�Z�H��qt*cY}�mr�\�47n�'�S1��@��`�,��H%�n=��{fTO�%6A��/g�ʹ�W1N�D����r��k[��Xp�����vKFl�r��{$*�|庌���A&b7�W����&� `������2L5���LBm~yeVT�;y�cD**�ieC6G���֝T�9����A'�l�R����gU�H�Ȣy�4k_�:
�V�׋���p�
�aLp�śr��-��6��� <��x<��R3g;�/��p�Ƣa��-j̩�Bx�:̽���Jcc�L�6MJ+�e���2uR�Sׂ/2���6�j��Ue�U���L6.{L�ɼ|t�||�������owH�pKg��Z�N�.�$8%�h�u����,[�@*�b0cYSe<2���X���-]�7�T���@�1x�I�����H�X&ů&�9��X��c
��o�QVt�-'������:{�ƭvY4�Y�X��LE��Rm*e��g��'5�ϙ�Oɔ��t�[�]���!v1��j�,�~����N]<[��ҍ��6�xr,jH3�i��2��I*K����Lb0�t���{b4.ׯ^���,=��
��>�[4�"��P�V����+*Vv�e�Z�G-��͊KqY�e;)�vx<��^��֕���8~�X��-
�l�1]�_$3�̖ںz)[0_�Κ�,���.�/\���OKՔٺv�<�i�\�v[�8'>�V�O�OyR�e���s}���*+E��r9t���=��|�OACl�V�r�XrLr�rnE�O���%�!3�x����sf֐��
����)�d������;:ɴc:��r��֧1!�p_:�S/%�՚�IjP4��)��P��B2�LB�$%ZR*U��r�V����ץ��OJ*&�"�(
b<Li(�b����(�`&Ä8͍k�{��Y�|�4Ϙ&%`�*�H��
�"����]r���h�)IL��{0�4cU�%2�)ͷ,��łp�a��	�	^�X��ьSC���egS����OB0/A��ڒ��Q�s!1�F3x��9y������T��dM2k�<�9{�̞=[�7Ɍ��%Mt��y�}���/S��d�W��>�U�;����t�h��x�F�l��ةtխ8h2#�J0gE=ֈ��ƻR\\,�yb�����l�5s	X�gչb�o�q��Ln`�Q~��#y�/��_�Z�������$��S��$D�m����P��4�4� 7R䭴���a���x��ǥ�!&��^���Oj�
�8��]��.�^��.����r��	�/&�5����!g�Tq$�Y2��OC�ĢY�|�<�y�4N���1��83�;��gOa�J��s��F*)�JUqz�L���H�Dz#�3<0�Y�\�K3��O���ʔ,�f����T�z�Ձ���f�ʀ9��2��Z�Xq��0��e �*I�����r��qe
y��-�p�|i�͵q�䰀o��n�ɑݭR;�Q���&y�彃G�㓭�d�5��gi�a���$U�v�K]e�4�^ 7Z�ȷ_������'�iS��:u�\i��N-E ���,1�Ҥ��֛o�~���1�E(#R�^-�Q�
6����s`yX�@dA��s��T�����S���[������%sen�4��0Dn�0�K�w?�a)�����!&/�O�k9|⬄��RZ^#��I�d^��
&��8!�#}�/!ٺq�l\�RZ���Ȕ�Z����>yR^��~9r������S�V7I�����/tG��]����l#�;�mV@`�r���Y0=O�z��3ؗ��F��,�&Å�R�����w:&�t��_Ĭ��a,�(�s�a���4�C������FV,[*7��9�gd�`������ȡ�ޔ�I�ԖU�i�r9yᒼ��{r1�'�<� p�0M�>-�CR���m;=,��;?�3'O��yR�Cw�b]8ccc�Ҳ�8�pR>>zN^}�-ٻw�t��I�|
�T��<�<8Ņd�@ؑ+��7�Aﶊ9�+3�r0sn͸�yxY�d�����/@��d-�dŲER[?E���hH���.Vu{{�||x����^���#42\��M@���0�ĕ�xo�W*b!ٰy�,[8[�.�#���9���}�˫�yYn^���&��p�,���XJRR�XP��n� V�S� 2����i��������42��+E=N@�v�/SZ^��DO?^wL�߫�@�/�������,?�Ɵe��e|@c�51.{w����sf���ҥK�f{3�{{�?y^���+im]�@V�o�_��B��\���͠��b���w&?,� ����g���L����5��8�V�`�n��k7nʅ��vX`�f�%�4��gaeAo�J��b�O�@0�7e����fO����*`9��sB��
h�~���y9�zN�~o��F��s�5�z�u�\���=L��JxE�2bLĐD"�Ca��9��!+ΐ��Zd��F��.��*5�p�����+���k�$6��N*J�4����@�i���F��Q��(c�7B.*�ջ"a�[Zf�ޙ4i���AQ��V�������
���18�����ޞns���G�%���0k}ii��TVA5����V�`|&f�'ʄgO���dM-Ͳb�jY�v�L�ڀ��r��m9{����,Z�X��?�)���ۻ?��g�a�d$a�%��n���3�@q<����Sr��%9�z�/-1H	���$���P0�9��&�B�A"@_[�`'�a��M�hT>5�l���XpU����l 5�L�&c-إs,$銠@���w�_� v/���{T�3��<��}��>X�a���ȝL��^f̐���Ʃ�d������e2�*/�C P���[�����ƕk�M�Ҁ�r[&a$>)�U���S0F6��~%a~H�)��r��3g�ܹse������u��z��8�M�����4����qj�㨼�\*j=2{�2'���3�'�4>��ڶ[7�����5�0��a��e��`H4��F�@gй��C.]�����߱�1il� VKm����/| 7�^�%k������P����r�Z��)Ї���
�\�#����j����C�����cOä� hU�s��{�%�Sq��"�e(­�2����?�cym�Guh��sgw
W'i�	Z����O�ǌ�EJ�"`���3��՞���)�F����y�f��Jt����a@!rCY�b�<�c�4O�&L�+���K���K�ͫ��Jej�$o0��,�r��.1=#:ɱ��$��bp��<���Ol\|u�/����!�:$��8�+���E�� ��Q0��j&��h\t5Yqԉk�N�*S��X�������ȫW�Jww�� ��A@�M�$�X��QI� �]mm���{��y��g���-��:��='�/�?zO�L�.-_(�[��O_yWv�?*)�2#V*#ɬ[����76��Gb�1B����kԕ�~Q	�� '�D�{����Fwʕ@>*�3��W�|�)��^'+�=~���N�Q�p�H�V&�q-Ɲ8Ь���H�k"r��>���Q͓J�� ����`���D}0e���ò�B����0����!)���IS�z5q�d �d��`$�����e�0����seŚ��l�J)��ae�h2!c L���:qKxh�� 5y ��.�!�L\���ѷ ��!$ �k��1}#��y<gL:֝J�0KW��(��4w�L�5�q �����k�/ޏ&5>:��Ή�ue`�����zz�@ʃo���y�-r��)9z�0�F�,\�Q��'dL�O_~">E��	h`{,�9�d��5�����F��A�!,���U�R	E�:���K��RkĞ�TB�{�Ȼee�P@ѥ���e~�% B�2��Z�R��e�4�jFw��L�d�J�x1��ye颹�c�f��1�¤��<�/ˮ7�R 754B��ha�ϫ,�B�0Q��� L���n�4��<��!�p�GaZ�:��u/ldUa`TW�OTt�������4xf���J#�ЀZu�5��k��v:'�u�b5�5���z��UUV;���Y���V,�������w8k�ri�=z-�ʸzE��2�,��ݚOe|������=�x������2c�)����w��Y�l�<�u�4O���m9p�ֹ�Q�mI�	=�@ ��`9r@4
S��L+ٓ�lHޓ�2�|.��ae�V>a�#mf�o
\ZVm�;��0ә%��[>�
�9��-��o��h��iV?��L� <ff����fʣ;6Ird@:�^�J��[e��Oꪪ@�ͺ,�JO�b�%���d��������U�+�V�mx5�����%
� ���o���K�J�u0Y{{;�S���Ւը5��G�����QS�	cuS�ϛ7G�g͔��3�C-))�
 �_4��dJ�MR�q<	��/��bp@�M�"�0��5U2�c��^��E�T"�}�{��.݄��F��x�7 �My��_��Z�H�(�g�I?��`�*�����4�v@~��[�"��%Je�2������N���H�ȋ��X9�nF���,V���ӼB���d�ޓ�ts�m߳��9M�9d��"����Gw-���)o諊Ryh�:Y�r	��2V���1��pMN'O��a�nŦ��D�i����TBݔɲy����m*�����G:4�e�������DvtuˡC��Ƶ�:q��,<��z����2S�&�)���NuwvS���Sg���Bh�"������?���<8
4�E�] �n��F��#�.\и٤�u���T�544��@\ٳ��O�OQ���)?������#�>�E��p�z�W 菜8.���2w���S��b�宣w\��%����}��PL��F^�[����;��x&N�)�t6r،����0拾i�>T�����*=�Pj�.��<�25@�3 Ąg5�+�eQy���K%���ӧ$12$]�7���l@P0uTЃ�,F��`�1��*��-��m�<���ڕ�j^� (����VY�����W�>�9�����ˣ����eʔ)�.�{ ��L�U�g�y�$Z7�2a���$VR� )-)W�2<8��μ"��nܸ��mj%���<xP��٣!����Qf͚%S!�S8n)|WT���7�����
�F���{�;wN��LnS�����������c�ත u���>rDΞ:����EгQy�_����b���A�B�pKwC{�F˭��h�����lg'��/���p�}�'[8,�川���-�7
�� +l3w�M��- �Z>��T����A�q����4Y>���� &�<�R
�	����*-é��fHzb>VtB��J ������O>)5��ȭ��:�x�Mm UI�}GVy��W��7ߔ��[���[�N���� ˗/W�H��>�Db\��S߰*�c^����¤��\�azG��8��Q.�!|���fa�AM2���M��P\�F�8p@~�W���7�ʕ+(NLl ���9���.�[YE�ԡ]��XW�\���d�}/�^�|��w�zGj��d΢yR[U)۶m�#����ba�ɪ�k$�ͯȏ~��n�a��Gʐ��@�&�-g����҃��R8��p���N}�է�t|Ή��ݛ>'�m`4���-�04f�^����N*��\
t�2U���s��7��A"���T1	�ך-np�4���y&�G�eJ�4ٺ�QY�t��%���wwɵ�u�9��0�4W�oޔ�����>��i�&y���e��E:����99{��$�O��hP�144��optP=..��0���e�g!-������FX@�kfW�de�<gH§�ϣYc{yMڵk������6oެg_�`2S�v�3e�Y���˗ɔ���^70^�̓�И������w�I6n�"�@��d�@NFn\>/�ф����T�����/�DN]hӴT��k��U8=��h�Q@�6��S���=��ҍ&�my�=.�w��/۲&���Xa˝�&��;�$�g�ɩ�vv�d%���e�̩��3��h���`��Ɔ%�h����X/5<0�l�`^����R��-�7����$w�|�E9v����5j�=����o˫����jɲ����������"[\�z}���p��L��̩j������ؔE���bQ��PQK�c�ڥ|&���F�z��Ì��U
��#rNH��V9�%�J�?�Sp�s����o�*����]�^�,\�^'��AI��6�$��
)��~�C�Q��E�v K����^u����6��N6��)p\�\�)�{_�>�I��G��,��\�эE�ˤ��ޫ�n�p,����3���tcy,ӆ�3�|��Ŀ��QX�	*��\N]������@�",�����Y�S�3�o��p�����X�u5���%�	c�S|�O#���%Zv��'��kW�[�jP� (� �����:��M-�}�k���/�6L"��W_�C5y���X{����V���:��2E���'S�e�<V4�hњ���:逓P���A �5VW\ ���G���^c| .Y�W�ȟ�Ęn$�@�'%vj����U�84���?�&�ر��v{���R]U�&���n�F@����b�^܄>���c��ڗ|�1������Z|����Нu��m���[r��	��R��_V^z�]�u�X�&`�8��9��r6]xL�0���2"�d������}���z�p8�Ӕ�{c.�g�+
���O�0���H��|�$7~�W�̰,�;C>��C��]���:jjm�X��`E�@ƴ�.�Y�+�*�LX�b��m�<~���j��_�Pc?G����gX��e(����H��&лb�7Ex1�(�s"��ėCx�%�r+����\����>x�f�j�TF&O���H���8�_J�M�!�ML4�1��5��x:���(}^ϙ"[���~j�}>5�=M"M�֒�����c�o��o�T5j"�Y����LֽO�~R-�IRR^&~P>:pZ�T%Agg����}���
z�!8@����X�?��;��o���C��;����*�F0���|�e�\p��*������p�F6��?c�4u�����I*���!螬{��s�LJ����b�)Xj�`P�m�Ƕm��������R�N35��J��Z��n���x"��.�d��� �M3�ҵ��{�0�����Bh�1����N.�����~�O�q�4I�~ǰj	$l!��~p2���O&�Y�ζs��\r&���J'�b��3��+��!��x=�q�}� 	,����z�],�9uXNZ�r�6e�$h�.M��1Y{��3\A`�!houu�>� ���,ӐE���[oɲe˔�y�+M.��� x���̙�9�U� `k�̩Ӛk���"��ʱ#G5 ������x���g%�d޲���<�1�ˮ}� ����r��t�����B��'+:gpj~5�
��^!y�pЙ��M�N����q �Z�H�1��X���y�h�Iƻ��%��a)��(� ���Q���2`��lK�qh*�x�)�,��>�����T/S&O�}{ߗ���F��o~S�_�)z�<��O�vhj"XyV�ÄRw��������~h��.�/�dB������GG���d�2)��"�a8�9ܻ����	X���֡AФ���R���{e����N�j���s8�R	|j��{�T�Aǀ���P�Ift�r�Yq���r��)yj�NGˁ	*a����-�%����&�EN=�,��;�7��n�csM��Ro\�:)�)"���Z� ��&��+2�+c��#1Ǣ�݃���ι���OT}J�=������q�>Xǳ�=v=���F�d���*$�Ӭ�:yf'��h��y�u�H[��`�2s�ԤqQ�(�l�9*.
�'RU_�/%�p�h��ܤ����ݻ!v������$1:��jj�X��#��k�{���=I=1��o�&_��W��o�o���� ��s��{�B�w�F�y�M.b�g͙-7< ���۷����왳���S"�<��,�>�k~�<j�z�\�pN�S�M��
�P�����,�2rJrh�	4V:p\.�bNk���h�f�k�56w�<Y�b�����@�6���8V*�3�����xV o�g/��L�1C���/�<`0��=�\l#��KK��2��/�z�e��7%xFڙ�@���S�a��F���X~0�B���)�v�[�u��s����舮���"IvHȓ��>�]r���|�W�m����&���[�X%�U6TW6���E�+,&��{%Z��˗*���?�(��Ȭ�-�o|S����W�`&�U��Qn�.����~�&�AcJ���d�i�̙2�z��)��� �)�G����9L�]�4���m�o�٧��C�����i'�FSC�8 '�Z$7o^;t�㛧�j��]zݢ�Kd���'�X��pH�5w�h\D�IM9ޫF�SxN�5��g�n�t�<��h�_�8L.߼~K����Y'��K�[���J��ʵ �y9t�yt�cZ�r��8��KEi��Y���Q��O_�s+�0y�p�{uǵ�0�n�#���چ�)�~���-P\�'�B`��'#��q��ϧ����7/���/����{wi�}II�ݯB�b��q*�*A�rGK1D4C���P+z@e�f:��aa׮]Z��g��;v�d����@��4�I����z�Çɶm�(�;A5M��ŋ��\�xA:��d����.z`dA��$LoW�m��fih���CnƝ9k����Hgw�:K!���:��:�X�H��?�s��g��y��i'̚�"�=�ƛ��a)�XD��/���Au6��k58Kf�3^164��"Мj��&��INoh�tҷ��my�?�2"� �q��\%�%���3��c`�bY4o�V��z��,��ŋ�HQY9L;��Ј���<�������V�m��O~-9���Ĝ�tݗ�����<�ܫ;�?���k���"��N�xE�q�D�ua�p����w�����4�Vv]p�[�Jl��Ih 4M-�qvVsC�K����������Oz�B�E�h���r��Qپm�<��C
�����ghhP�C��;wV���lܰN��͒%K`c��.�k�Z��?�U����QX�4�|�<yR�6��=��}G��Q��߀�IB�'�p���D���<'���G�M"�fƌFeI�?nx%�VVTc�o����|�ݏX�AW����R�{F�<��%=,��"(0�v/����/H�:��Dc��ɝU%`ݹ��F��WV�$y�?HKe΂%��0CwDs�Ξ8"�0F/<�CN`a����RZ�"� �g�2ܝ���3�|�Y����ex��mi��=�����n� '1)�=�Gd(éY<g:<��r��n9��~i�4Ej�q�g��zθ~	Ot��s���X�W)���q����i�l��g�\�rU����d����	�Cs�X���F������s�x�y����_�9����ի��`�嚵�tcjoo���CFGG�j�l.z��p���;^L����i7�W���@xr�Sr��-ux�Ȍ�&e*2* @�'�"���K�9{�L�4U._��)�M-�b�*9�}�(�[��<�Q(����;&��N�D��LJ�2�������J��o�o�����J�uau��� �nܸIn���SWUV�B˙���\�5|2f�����ɡ��e7�P�`�-��E�)׺��g�<a�q9�.�x�30֧��|"gx��L̳���F����Ev4��H��c��i���wJ��˲�פ�_����Z����0�O����SX�Sc2i�4���ń�́��0�̉{쉧d˖-��)p��w��V �Nk��c�Ɍ��r��Yi����D����$���/X8O�F���羨ڌ�������������x��L�a(��{�ͮ��'�B�p��j����,� 0����ʪ��v�`�iZ��Gv<!M-3��kr��E5���^�d^C4L1���-�=�3�n̳F�`�����߿�����_0��Mo�G,�����+�]��Mҡa,������Bbhk��q¥�(�۷[�����������rk�M�j�l�L��sL����BO����x�d޴<���0�$��p��q���I��������e12��I�?&�K<!�Ei� 1H�^V�B���jAx�#,y�M�{�SI���>�l_x�9��E�@�X`,�P��ӧO����er]���;/�7m�}�gr��G��C[�u��S�<��#:�<���f�����:�Q+t"��і�Z�2<2� ��'��zF�f`��(X6�vMmh��=L�wt��-��E��g�\� +u�ǇNH}����ޞ��z��.+W���Vˁ�wˇ~�y�Z\SQ^���'NSFk� oO_�{~�W����?���t�?��|��_�~�lr�p,��1F�������o���m�t�"���q뺎��G�b�-3푥0�5e��s�v)��?{N~��	I%Rn�K+i8�Fy�8Ҷ>X��~�S&��r�Xj�h[i� ~�κUKe��{o�,}�-�Ӡ���r6�[����5���l�h:��� '�4 �U�SQLS�r�f39HN2�:m2�w;��EM�ѣG����?�U��}|�j��M0k=rZ���_��N,+'֭ݠ�cY��KW���ը)y���r�f����'�}��K�c�C7�4ˍ������;'y8��Ʃ�jҘ������� K���!@�>�]�c������A�oٴ�|H��b� ���2wYVA3��ʁ�x����w��]��?�se-�z�X����� ���7����jJ��p��G}$���JS�\������fA���gd}]�<��Cr�J������˩�@��ѭe!��O9m��ɏLӼ����Fڳ��)4-�%!y���r��Y�:�Z]�^.���w6^X�@��?��CS���b �i�N~q�8�o۪�e�˭-'��� ,9�9�Y�%k����Q�^�N�`���۶cB����ǎhU@��կ^V3I�@�f��]���2�e+Vha ��xh�c�o~���X�Q'�ډ��[��x�>>�pX��Ύ>9�2\t��m7�7�y�x���6�=��p?@�Z���������E�N���3g�9�����ڞP��\Ȯ<Z();w��}�{����<e�� D�+�*��Vȩ�'t��Ff8��o�~G{<�:S3�����[�lA��_�\:�H��8T��5k���s���)ۿ|�`��82S��)��?�*)���N�d��ӏ����W%e0k%1��ΏT	�,w�C@��9K�	1��=��4�}��)��~p�
qN7��B����*��z�ԩS�]]�����CKq�a:o^�.�O���*��ۺu�Nd*���_��5x��U� ����ղ�.���V{�n�d �L:��Obe�pg��2?��;��ͬ-Ro��v����DNSP�1�S��a`ltX�ҏ�'8�Ɇ�K �1y饟@���g��v|R>x��V��kf�z��`,'����XT=m�;�����[���T¬�>�ϟנ�m�(wKaQ���ޮ����<�ڕ���p�W=Ϟ�Ae���yh�*=e�ąv��yF�2�A �D�#=<�������{L3�/%]�,��#��e���{�_In{ä)�@dz��b����uOa7������7VVQ���9,c#�d���*��#�����U��X�L�y�*<|��N��(��͙��A��O�{�\�"Yh�nx��p����4��=f��u꼩ST3�7
�Y�b�Ǝ�x�'ZѮ[� x�)7�c><���@S�Z/������auX"�Wo^��[����R�������ݡ��	���!����?�6h�����<�Y�[�����AJ�XٻiF�f&~���I昰��EQ;
�:��ճ?��T;������|̜��<]*��`g�y,�+�^ ������oɑ37��1v��a���O;�/z2݋��@yD����6�%�˚��$|��!���ʸA�Q�LVc1����&g�wtN����$/�S�t+�&\�k6h���*#rRi����J���8�,j#k�>}
�>�i	F�yB��%���G2ٔ�<u\�6k�e���i�Ih��,�@�P�/�*+Q��S��tH� 
'���K7�2py��P�\���CM�ls���9��mܸVOջq�&��zxW�^SʅA���A=d�[��S��`�-��cj�.`���[[��@\V.[��T/]j�����0Ŵ�տ��n�|�0��h(�{JL�0m*�����P8a�oܺ�����Z�|������dw���>ؿGvV>�>��T�Aێ�R( ��,����r��u�r�*�8��;�����	���|���ADX9h��̞3]6�[-���we��[Ι)�,��	��w���<
�HQL���c-�� 55Ks����Y�Y��'�qձM�b� 5Kv^W���I*Hׯ_/_���r��Yy��Tl�|��������YU�p���u�`�9sg�e2�?��e���Y�Zb�ܙ
ԓǏ�e�-�����aBZ%���X��ۗ�����̼%�o�z5*�~��3𜖲�IRYӣ+��Y�ɋɕ�וm��kߐ�J9��樹i�J:}X�d<���!�<y��O���\���Z5�ƾ'HK�B�ˍ7k���ŪeKefs�ik�%���(37C���1�p�.�^+ϕ�͓��q����+�ь���pC�k�]�P8g�`��`�>��<�c�t޼���[�HuY��l�U�GL�D*�6�c��=���|N6F6��0<�V;�V͕��|Vk�8 �U�+�� �B\�۶mS�E�x�b�i2{0��3gjUg�j��4; r������\���Y0~����7���q,�K������Qj��0i�p4N���sa��	���O�eKf�¹�x�6��m�vwu�j]%DEy���X�y��i�j+�c,!x��/�gԴ4��z�={��B�/^RsG��ѡZ������3�~V#��~W�\%�pȴ��x	�?��?�������_~���Z��� s�dֺ�S䩧wʋ�����X�D����M-��a"�O�TK�\>{RVm�"�V.����Ϙ��Q?��޿�=�Da��2�T<��V��퐇6���S�����������Me��Bݏ&�$�A�:c#�p�k@�\Qd6����L�ʒ�Xt�˝��\^Wh�' B��v�4Ή�] }�Ӵ,�|V�~	��`߼y[���Zؽ��o�Q��u~Q�Q;�Z�ʩ��SB��k���|֤Iu��;WY���M����E1�7���Qh�~�/����)f@�i\�C��khz(�zu ���Fܗ¬�̅8��X0k���3 =~�~��;o�+O?��^��/e߾��}M*+�5��� ���Ď��R�N�������9���㢛l��d���n�zy�׿���I��i�L,��I���4��.�To���D��[`@���<۶������c��L� ��I�J�k����-<�Ա�2��N�!��Vz���	\�՛3l��!d�_O��Y��!c ���h�&pxs���эk7�\F⹺�zH���>����,'9q�\�~S�'�&�k1p�7�˓O���|��G2���Uٷ�=�Gb|��P3�UJS�f�:Y�z��>sR._<&�)�oQU`�6c����F���.�1�E�<�]�KW������V׫���C�u�t<�=�T�Ν�s.PM�c�Jb��k
�'��>Hz�4o�V���?�+ׯ���ɍ����l��.���2�?���,��SOh�_|�E��;Z��붔B�`�>�ltA��XX�P�`�Y���Z���լ��0Xs���0.��s`�t�$��b�X�Ga�-����<��U��v�\�TU.?���$�Q�U��^�F�ǈxu�cBC�܁!)k�@��ժ�X�Iώ��19��427F3J3H��ǔ�=(�Ϝ9��Aa�� ��Z�=���S��O7���C�0sL��X���y�=۷n� �Pv|�G���J?j��g����t�^����$����l��G&�fS��g�q�)%�.��%���J���W+�,^�{�\��[��A](]Ъ}C}2o�"=��E��|�YOd�e�Χ�y��~W|l4!����2 Ǘr�It�${���M@}��/�ح`��[f#8����)�d�C�!�T�-�-�ˋfHoW�m�fCN?*KVm�c�@�>	�3$i��r9�]�c�'����h!���7����[�ƕ�RW��8�l�p�p{C� rg�a�05��$Ro�M�-[!kW���헤�Qe�D0K�����j��`+N8��SUz{�5��z�A���	��ߏ�@8+C �:���5+��P�kW�ܙ����z��������"5\�4�'btlX�l٤�g`�_O�Y�z����x�U�w���2�e!LiX.�;�W
V^�&���Tz =�1/�������~�|xDZ/����<��4�E{����+uq�����������W^Q��A��;g�,'�	��;.@�����?�O~�Y�f�n4OfT�U�w��B3zύ)�]�n4J
ښ�446(8��s�Γ>:���_�D�΂��KJG���/��Sg�O��$h�����n�J%���*e��&����R�Z��g�pC�Wo��AV ��Q��cHʫ�lܼ�s��i܇>D �i�u���ZQ	7�Bf��$+q�h�!��Yx�Cfc���8����L�2YY���Y��0*O�����ܗk�:w����Y�J���rL����j	�\_�Sr���Z63{^��>w	��M�7oި&���C��z��'tw�0*u��;������Cr��yY�n�TW��M�tA9{���,@dYم��G�m߾}���b�\��}�/��'(X��ki�f�b����ߪ�?�zQ��e�bX��Y�k�ya�ǜ3eJ�t��`��+g[˼%z�٩SץK?J���|qoa����DЯ��E9;#����k6I|�[.�=!�E=|��q2�Φ�(���*�P�PH�� �$�6UW?I;La��h*+��G�y��\h&(�*���X�u���~�3�
$ขɠ�lj�y���s�,��q�����8������?^�b���dep�/�?'.^�Lw/�>	���niiV�̖N����;�i�ݴ����>�%M��,����,\Z�%+�!t��	-f??:��S!��
�^cbT����ΝՒe�dX��mø�g��K����l�������e��i�߼��'��%G�={���e���	��0��J_��Q����X����h����q��
���
���!8����94\:���)�3���F�X�� �I0���elf�t�u�25����^`|Y~*K(�Ӓ�(<��˗��㇡�F��,��#�y��׭[�G��350��#�=��<�{σ�{':@, @���FSՒ-K�c[�؎s=���N��;��{wfss7�ؙ��8.�*E���;�J���^��΋����#���}��9�9���'&֊�0� �T()!���i`�J<���w0{S�yPTP_���NNN�f�c�H���sg?g��[x�
I�. 帥e�v_#��`d��iV��HQa����HDX��<}�\�x��%Ղ�%�����?6m��(�cS*T�~JU0g%'gA*��*�^��شE�nH�>˰`� �m�v�`�޽�H�T0�.�_\���n���,+U�^�~��<h�+~p��b`�Au��V��;wU�4����,�Y���R�S���^6�d9���e<�Nl�¾�%��:��V�����8033�beˊ�1�๡'�J�����+Muu�]��}�yr��%��s������7���O�\����5����[$N1ï�KX@���`�&e�тޘ_H��z�IS�Z�}���O.΅x��������61>i���P|UR�px�Y3A�j��X?~Ҫ+!^�$[Ɇb7Z�&Ƙ*1�#O?sƜ��|h�s�N���3��cB5�w�XJ��e��얙�U5��?t�e�O�)��ƛ_Vs:%]��9�o|��DGg��Q̱���8U�;�t���	=dQ�ڛ�ScS�\�,�K�V�&%�n��kT!
�kū��Ckn~P��YV�	u��}�yz;��/�������0��sE<.%9��Vn���P��P�������?�O���J��O{>��[u�aoƣ\X\�ֶNٞ��CpT�H�,{ftBf��$7-J2�Bep`R�ܴ�g
ւ��Y*@���=$�rrd\O`�jX�@�9����9=��(����W$l!�[�'VB�*.!�N�c�G��uu�1::fm��vXw��ꢕ�t�&��'��i�P�2��W:���ɁN�8&)
,��S3�«?�����U�ٲu��������V��k�z�v����?P�Ԭ�i2/4�/��L�t��ę����j�P$��_��Lě�v�H�>֕L9Oپm�uWW�6�oi5=���G��:Hy�sP�+(n��̅�9���4���C���$�R���'cX�zU�~i� �X��P�J�#�ѵ�ղg��U^=q�>C��;Znb�
�T�_����� ��*�C�M�M��@�j�¢|)ؖ��������g
$ӊ�<�����KTu�s2Sׇ9ӱ���b雅�1'F3�6�М��a\�\�����9'��M[˓b4j����!ج��߫�䱣��,?W��$�;M�~���O?�ؼ�T=�9��296��"�IO?sLMT�ܹ]"1�q�W����{�T(&�h��e�����6��>��k�&_O�T�?T��O���c�M��4+��6����"�mMV&�	�x�]�.�x�F�(a�c���Ȗ����(�N�#��(����!�R��7�7����hK}5��&�>����\����nx�\�xI���ckν=��)�"X�UL��(�$�����7��c��p����YN���uu�#�<4z��
D�V�F������H����07����������1��~�zq����d�`�~/��D
 <Bh�p5iF߈�T�S������RO!��0eOG���{*+)U`bf�_�cow��m��v�کf����S�Nȼ>tkS�4�7������r���z��ګ_�SK�BUX�[�6n���Jբ��R'�Y/++��6#��ޞ*�}��ӯ�n���!՜���*`3��ZI
�}�w�ޗ�� ٹc�E�kjjU��%{�yz�/]��.R-M�һ������J}�j������83�`�bl|�j�'PG�\,��h@pI��-g�ļ�^�����P;� � �Ú�S	{ི/hg�yguS�R�y7a�w���޸1�,@�Z3(�w��0�+N��x���`>C�V������B�VЎ��Ӆ�����J����1�M���|�4��' ]o���؄�L89�x��7C,���m13;g��Bv=l|
4��MK��#N����V�¿�� �p�}���!�U27<���a�R�`h��{Ŷ�!�զ�g�P�N?E�n�X��
��$*2ش�L�_|Ӟ�̌j���
epH�j?��������F�QFN�fc���u��hT��@�T��(K�*%y�%|�#�%ng����C�ol�g�)Ǐ���6���"�������K��}���������6e�PB�$(h*��4�!�UCs�KS��r���fAx?�~>��'����!%B8M�2�epY
.ccb�gg�>S���=<��Q��fۖ�Rv���4��Ӭ���'�4�
�d��0+���b� �e��������1�D�vI��/�,�`���nIV��*�Nd�U�f'UR��J\,����!V�g�zz��(�T7�����.��q21=�'2�b5�w�.���a��i�|��*H\L�a 6���(]�����s=�m�҇���,��/�;���P���͛��3�JC}�����L�UhYJ��n�n�kTl��<�uIO͐��eR\��4xlܼܼuG�VY��Ɯl�{��y�$�A'���4�����J�v� `��m��C��2�=^��yľ64�I�:Ad
�y��b�9-Z'ŇtY�1��X/{�-������}�����^���ZMPU�\S��Y�A��J7��y.6�I��O`
�c#�}���V�bQ�)��4 (���i�RAD�"`�۬���7Cs毳�S�V��#�v]#""�����K���W_W�h�WmjRs���`��K���C�P�z��U�<�f��,�<4��55Q�
G\�p�8
>��+\��� =@���[7���l�oH��ܻ{S1M���}�,�G�v�����R�T	C�v* �TMVe�[�쐣G�Hգj;\gξdvL �V��o���"��@D+^��@���,�t��t�w�frB��]�.y_��>N,DNn���Rm�C��,�amF�3`�ٖ��:�Y���rtq����DJ҆.����r�?i��ڤ��T.����)#���XR���� �)�b�l {H=B��< i���fiQ3���nf�NU,�c�;�TC�0��v:b����ba�v�Mjm��D[��6�z�`T\��u�Q*r�@Ϟ=c$�/|��뼜>yԙ��'����I3��>��������%7Fi0�,�=՘��)z��֍�go��RX_?���Q+.�g���^M�&9~r�j�!�ܣ!`d;b[�{N���}�T�w����p��Pp\n�,!q�
O��X�I�����!b�R�KYsë������>�����w��-�G��۽��>.B���,��a�Kf�o k���e�]k�S-�6>6:ر�
�L��ᱸ�����p��) Q���}�����J��q08�v�jRƜi�b$�xF`��5������uN<�P��� w;7����	�B+?yL��X�w��i+N^����7�YZ\�׾�50)$���jTLF���@j�����z�a�sXd`_��P��gO��@�b7oʳ2�l��C��f���	a#"������������8�Nii�S�mVf��֫i&��s�e�Z:�"�MT�j���r*'��urt��U;��΢B	���x$s�Ӓ��jm�s�z_���H�hk���G�ɘxʙ1_����G5р9OT����~F�XW�ͥ''��z�$�������Ң���dY9r���[�4&oذ�#����|���&�v�%o��8�jXb����=�!%��,�/d��iǬ����k<�k�9,6Z(5)�6��Q�z�V�5��<�|��5q<w���_�)��m�M��ٙy���D�P���1ņ� �g�:��s��׾�ا��8�]����lU��h2po��KE�#1Pie���逸Oii�ӜT�ܭ��/+Cr��B��Z53F�q��.u��ԅ��)r������G�̽�	�����e�Kl6��A8:C��P7)Q၊��lD/�ވ����w���V�0hHO��y~p����XJ�*B��~��c�
y���� �m۶��=��o�N���c2��p����ޛ��;_�S6���<�V�?��_��A��v>��%=��/A(����ʧ�jJ���l��6�qK�Q�6Η8�ܬi:2�xFhT�.�s��PE����85-C�Ɛ�L��zESs�qnKw�������� SƆ%/'ע��#�ҩ�P�s��nB7nݖϿ�l�Q���Y�Q�>r܄ME�?�y�&�Y�,t�W��V�R�j�i�Б��Q�=�zF�qJ5/����6���2
���d�*�_��7�EH��8ʇگ?�F}���m^h�:W�{F(B�,{Y�[{[�\�vUv����>�F!���_�k�U�&d����ߐ(��Fr��W�3��!�������6��=x�)gr�YA]�=�<�D�ҍ_
����@q\���յ�+�5�d/gX5�������@��A%�"H�8�gh*�<Z��au�99��f^�y�mSݯ��-
L��}��3"����&&�R�|��uk������X2>-85���?�v�?��?K�o��:~��Z��� mIY�5S  q�I�����;~Ć?��8 ����2;4<V^���a���:$6tp��)�Q6�6�B`�{* �Q�G��!�Ox&Q���������=O�?gdp����R��KLl�u]/��DM�0�PŲ�6"�:o���M��I��e/�N�:�*8�_�Xh��%�:֜� Ȃ���r�"O,�Z��?�T���b}:�Mp�aq�:r 3����Є�W�b�F�
u�à��.��W������OZz���޷l٦B�AOH�M�@0)wƻ$7F�.*J^�̆zu�{%%5A�"C���L7�SOn�EKq�ʩ���eA�ǝ�j^��;�]u�7���R	�Tl�߄3W���L#��F���ڰ&����δ�I�i2:�� �L��/�����Q#Q|G�3��
��	�����RW�U��>Ňajz��3V|S�P��cپe�b�i�u�VC�ٻ]�ِ�=0���'O�֎V,Zl������7nUşT�b�yk@��mcd��E��
�!Rxz�r�sMI� h��i!#{�f#����746F�q�g
�^l>99���(���ZDͫ���%+Av8q���lEkѺ8���f�9ry�Y �9�����xhN	M���dN�C�z�h�i�hq��媭����KbT�Ғ�u��-�[�%���j���eZOnfZ���=~�%����mN.���}x�ٳ��=RS]��*e�6����˪$9�G1�!;\��m
�We��"�N�R�Zg@��K;��`6�4�{,��A����J�۔%���Q�쁕���.I�q&($�s�6[ܮA�驹E���^Y��&ʿ�կ˃��m��|�MsB����Yh��1x`�1N����a���3]��E4�z���}rilƣ
������N���t����o����j}T^����y|�S���a��z���-���6��$p�.:���`s�|�%��&y?�ƃ��V(�����^��Ʋ��A�d�����>u�~;�����H_�\��.}aZikQݭ8b�<�u$H���P��ܺ\��IyE�>�� ����
�<�����f�՞�.�Sa�)xfzA�V��_Ń��U��Ip��.z�01ff
N�$)ض�>��k�&�1�J��8��SM�Ei�}d�&35ٺwn߾/�)��6ԶI��ꐈh����ޡN������E�P�����J�5�y�j���b-9��;a͌�0a��C�}N�J_�V��������A�CxǼ����1ﶖ�-*`����]�R/g���O��.�E}��a�l�F�M��^�a�1hT*��iw�͉�9{
�i.u]v랅�ʒ���a���`I).ޢ"���  '/33��F{k���޷)�r�t�e�K�ñI��oHL���j�f��iLx��|K�c]�UI�H�Y��O~�+��z�x�7 TZ�;��٩�䞩ô��
�-P[��4@lT�
׼�F��Y9�����JU�}��3E�
��ާ&��/6��p�xW$ۛ�jl���������XP�vT�<����={�ڄZ����6��ד�m�{8r����Q�,��:7{�1b)�fY?�CNM�Z��u&�@�R*m�z�)Z$��`��B?:��!ƶcu�8ak��}D���U�ÿ�L��;п�,:*Ii���T���B~х�c:k�邶�kj�ٔE�b��-a�P��q�Sy�7!?`�`{�C]�$���e`5;8ԥ%����A�mb'〺�[�檶�k��g�>a^3�;T :�Cܶ�H���\�vO�Z�͛d:��^�W��W>��Փ^����_��K���-e�*�cr��)��UQQ��oB~؈eoݾnxtx̪3&�G*�&�0N�"��3D5�z��r-���/).3�H�޽=C�9w����iŗ7�\��.�s�� A���/�|��j�j�l��ajG&�AE��2N��"0�&!�Ev�M~��w�@d����(;y&�G,���uR�eD�R3��V��[�d�.Ft�(��1�S�w�t���᠌�Y^2M?=7�3����D��Y�_���\%�a�EPZ��KV�]�`=צ���Bs���>N=��U�z$�V.{0��fY��UՇ�ɱ�o0�R)�����ISÕ+�ʭ�7�����YF�=��K�v��#�9p��m	�����s���\ܱZ"B�K����AFGf$7g�̪&az�����Fݱ�TDǄ�k��j��S�z��d����~p�؞���$��Ԥ[�#5����Č����D*.��߯�ҡ�d�r��.��O�:)L���eppL:.G��?�`���g�<�䔕��H�qw�7�fJWG�	&���ޱ��uJ��a�bSd��p����`���y�.�,cm�O,��
�d��׽����gF����U+x./�>Q��g�W�V7^a�Nk��`��uB0����[g�����ͨpT*����7h�b�z��{�9����˲

j�;��R�w��Q)Q�sz��I�fyX^���8��b��Wo����F���@q���b�w�L�:�Z�ܢ����erb�4넞��=sL����bٽE;�����O��X�+����B�K+tѧ��6�GK��O�o�d8�xŋo~�-��\RZ%���ln��c�iji�U�e	��
���o���Yfv��}��cvY;	F����HFZ��h��{��m:����P����|�8��J�)��А���1�^-�,�Ɯ�ҩ��p�N�6r���x��.e�X�@���=��s��AO�ŕE5?�!Ak#;��L'py\����{��g�M�{4�D��&*�U�H�[�t��T^;~�0�
�_|Y���~	�-u񝝽V��J��M���t��I�*P�U����8���C�� �V<t�O��IJB�ܸ~�rh9�@�w5�v����Q��IOI��jhj�r��������+4^X5��O�E��d@	M���T�d�!=�|�����I�T�[��v540,{v�SO�HJ�������^�'w��G'GM��,�j�5!A���2���?�������ֽv�aN��I�Qb%K�<���}q�\�h�o!��7N�{e��~zm�����Ĝ�k��Z�����;��(�X���#kS�]���#dļ,%N�!������Z/`zV��OqY�C�
�$���\\|ג�t�lHH�ʲZ51C6c��p��G��q����b�ȼՈ�X�]�Խ�wԋK����&�^�٩'2\>������á��*y n�餿�	u���dڳ667�g��d��K��ҩ)��9r��i�Y�}�X���ʦ��ҤNU��i����IIy��רr�V,��;�Y���/ݦ޾N�PE��رI�iu�;���nl��`�O��¼Z}�z�[��u�,��hi��E*SkC:��-gV"�0���K����"
�wm�:��o~~s+��fP�������
���q-;e2�`y�M���y�n>�e��˘j�$W�H�z�Ƒp��$�����
��M,{�-�����3!,�_*mͽ��c�-��,V�T��+P�(��4�sϜ�ώ�[�n*�됄�G��^��v�����\#���ge�J�~V_o�t*@wI]S��TV��#{�Cd1��P{&N�����Vq'7n�W��h%�a+S���X�{P���7뇕����9Yyr��M+m~��/Z��������ɡûU��
�j:�+����بH��=|��4��G@�w��]+NMM�*Y�4C��Q�b`��,<������8�\�9<��s��b8������;�5�0��p�HU�>����M���~^�p듬\��J=�	w)'�k8�q`¦�ب���=c�ihe\	�B^�K�\@5I��ȰzkS���2$�����TlUutd�͡R�CL'##]N�8e!�{
�����ܻ�����cD���Ⱦb�������/K�: �M��h;|������f��_��
}����\rR6lD�j6��U5��������B��6��;*?��3�ǃ���Cd�m�S-աۨ�X?u�p���یp���ɘy�Ąx�ԃDF#**W�|��:��5r�݂K���A�3l�ߌg~My�8�P�����I3�����7N�����I��0;��0Gs'!�X�P��u/j=�0�xy�fF���y�������;�|�x+gS�uJb���bt#�:��[z�>�!Ȓ<����W^zYq̤�W\2����_��nL���K��qZ{��F#�u���Y�X}��QQ!jf�m �}�$<,J�K�ʹ���뒐�$��k��R\�(H[q��8��ɵ�er|�X����$3c�Z�:7��˲w�.		0MD_����jB����v_/������(��sg��DGȝ�7��ED�&à<<@�[ne(�yN4UcS�A sd:dCr�iC���S�h4�*�.W��I��!�hv�@�u��⽎09���^�y���g������n�*j1��]@�.[�~[c���t��iC�����,]LN*������\�I��׮^7����>gy��]�89t��.x�.�5�h�l`���)+}h#x7oΖ��J��o�ݜ��z��V�y��Usn��a�!HD6f3�2N��'���£��Q�<n���9��)]=�Ɯ�p��)3MS>�Ve@W�Ⴧ,����^��d㨮X^���~���P_�H���%\�kzb^�j���Y�B���}uM�u$�������}+.��"�g��sP��T{9�L�&�֖�r��I�,?w�#�;��m�5���u��z`Q��7`b���'c
��i�n��ɵ�z�r����ܓ�s�sY%pյ�ˋsh���Q�Vi���,�}��=�F�~�2qy�|�ӎ�iP��lS��by9T3�T��̤ʁ���sgN[����͙�nq7�����1�\���@��G����fuO�:fZ�EA��ܲ���)$�tP��o���T!�ХZ�@��i�h���f����P�"q>95o�<��8@����jٸ1]?sm���	zFj�
n��նH�:�*DM�-�����:%�)�Ⱥ2w���F�ojj�
r�E�[��Y(�iTt��;�c�+C������	��Z���{.��K�������-�s�*�K5��,��(X>�K�6�!���6�r&Hh����4Ϛy��
_�7C�x�W���M~�w��{ߒ,�R�)yTUc�9����^U��MDX������
e<�qa� z��uijl���Xc��H��W��sE�8`#HH,���w��頡��&
6���WM�e�,{�������b+�Q\e���]8.>�ʥkUHvV�=|@�zz��Vύ
�S�)��Xo��'��җʇ�2<�ok879#e��ef���Y��^�]5��׊�y�Ν3煱v�j��~)(ܥ&,��(��h�a�k7��3V˶(?���U�9&�o\�*Zl�@�1�8G==Sz��+65ֆ���c�
��ʨ,`2���(\E������䔎~�2YjW #@ܿ3�Fb����&�ka���T�뜐����j�H�k�+��G�j!0��{�ژJj��9ڔ�g���fu�~t��Q��s��O�?e�):[�<�EVuG�׃`ce��p0II�r��A3�,&ܞyz�A�r��}K����׭�	��g=vȞ��i��nG���`"�yx(�"��\/�c�*�L�����u9r�ezzdb|Z�b�?m����J���4��0e�Y�[��[�B��٫�H����J��0���{��q�~�0���-���8��Wg �����w��n�No�3���f��o�Rr��������.�{-y,<Y�T����u�;�"�)��]a��`*wL��NN�ߐ��Aڑ|#ZS��t��܍&@?��?�Q=��;!d�)	�J�Sw������=
�=�&�ώ�9h<uM
bW��ge��͖k;�����Mt)�3ǢSgD��o~d�ɱ���u�����i��FԘiy}׈�z��9	P���jʘ���̸����d���6ַX��G=Ӊ�9=���/\��^�QLKߠ���BF�����Z����;�ٻw�I���}l6O{g����m���W��6ȩ������6ZH<�v&�38$ {��˜ ����0�����1o.H��KK&L�#������x{��'k�%��[fo�XY�S��u���~7�z.����{8@���t�Z�)��b=lyE�����A��`aqF5�3���Njj�o/���XyXYk�F�IS�CP0Z[�(jn�C������G��R�H����V�6l�g�=c��^�a�^��Ss�e3��}�W_�v���+��ݔa����L�&�|76:N�CB%@�����+c�S�qp�K��I�:9��������[ZSy�yKR��Cz�,@�e^1ߕ�7T�w;��ަ͹~L|�4��$̱��b�>о���z��p5�p}��	��^-��k�_l���AӭE�:c��rq���8H8�g?-�J���⪾�����e��U�F\�"˽��x��=׾�A37q�&� >�辴��ø)�Ѽ���`��I[����֭;� /��y�R�O?6@Lu�Ǌ�+N!�G��X�)�W`vnQ����$<4J���[Y��_zU7l`����c�v�r�3F���R�&��Ǫ��ͯ�,�y��S��kO�%�����ZĚ[ddtLRӒ%sc��w�'wO�T���]P������n���zJ}[�L�e��!�6���w���TMD���m��Ϝ�,ŝ��F{	��V�ЈH�X�'��0u��wޓ?���,M�ƙ.�K�6}��B4?�=C0���)���o�	�G����k���4��*�sO,�pGǇ�'mC���Q���lj���ZX�h��n��R;zj"�ͣ!��`��S��5�+�Qf�͌�P����m�8z��\�芙կ|�������{�K<��Y��UO!������;
�[�3�n���k+���D��o�LS����놂� 9}�y�W�_1�My����)�&�1�֘��'J��GD�^��ۖ�ƬS% s��pF��~��k�Փ������1[�j���M
w�Ilb���+Vk���׊�~�_X�=�s�@��-,;������9ռ}V]����}��� !>ƚp��ض5O�V&Y�֋��$3KF�D���j)H]h6�.���i*�7�nq��Zc�[��V�>9�D�Z]]�
	���v��s*T6:l=eC.��%* s�S��ϑ�!�!�`�l��
[7����.IH��)�,3,�ܙW�5����my�dcf�e����$��HmC����'�"�M�o5�/��Y�����e�����/�ݏ���+2��|Ѷ�@��l��{��@xHRj�͉^Y��ڮԔxk[���Q�}���-�K���>z�Z��u��âͬa���Ԍ��F���.�u\�Y*�-].s�c2<�h+ƦF���5[�e�-��o�^��hQ��N�����]�~�����}V�ME+�Om��`����mpU���9u����Y�q��-�eи��ҭ>iS[����̇�	�.)�4��m���:&&�0(#�N�TR�䨨��@�V=�7$x4*�0����������ܤ��pcY�D��@��Zjnn�L%���4~����bPzÀW]Wm������Sj�JH���Ӟߥn��u���}����Sa�"�5R���x��f���|yTUii�<�&����7�)�m��ɮ�Vc���N���	�������t}c�K�j
�:{���j�`�j���B�աa1�7N�w�x�ƴ�/����3��Fs��!�(�`�W�kxP1*Igj�e��(!�W��f� �P�������FuC<n|̨U5�>²<�f��g���4� �����.�{�|�>����3��H�[֌����$����^	�	�.�Gp���=g���Y��b�P&�X�S�����s�9B賎�x�V�7��=
���Ύu`���.U���m����S���.Y�i�] :���lݜgC�jjJUK�D�Dʫ/���@����t.��|�v1��*�!/�.]V!��	`;�v��������:,�>Y5�5��_��쭺�u29�)�
�Cj&ib|TR�l�W�
�Z�	)VYUUm�HB\��K�z���@t�0���}���LH���ݻ�����q	�)�6�r�p�GGG��Z/=���e��ֆLe��ҫ��Xs/E�~Ϟ}��w3yk���",��P^<v7d��ͥ����{�bi^�&��7��}<I�TK�$�&+t����M�\R/S���Ç)E��v���o���\�!� n��m�@��X5)ĥ '�PA�;�p�3s�)O?s�Nǃ{�̳av!����"'*CO��������w�p�#�oU�3�?%;vK�
c���X��W���d�맶M��mڔ%�^��''g%ZM_�:?��U*��Fʨn<x˼܄h�[__�����@9a�٢f���=�0�GZ]]e��	q�i��Y��op@i^=�!�oDs�:M_ a����3بBA6����i�c׮]���6���Wե.��8���k��q�8�0ߨ��n��^^�sZ�T!����Yn4yG�1���ȨAńO���Ű���PT�[�@?!�^�	�3���&�M����̉�����a��`��K:�?�"@8%�I�)�9[�CKJ� u�5�� bq������:�t����I�2o�RiZ�YH�
l��}&�T<ܹuM��@�L�	hDrb�x��ʏ~�+
�ԓ�=`�[Z�2@~|�1��F%�dYy�v��_���[��c�y4j
󁖌�U�WzWπ=�ᢝ�v�ү��07*i�	�r"�~��5�޴I=�g���!�;��-j�X7f,B���3uL��uG��)7���QoF��T����+�g��U�*^���2��a�t7;�7Be|�k������	s�TPaʆU���g.*"��D������0�.�� ���Ǵ���y�FI�bF��f�ٜ����%�b�*X���YD�֐*��]������0%����)HG��W���uf6�Y�k�zX��9��Y����oZlqq�b	O9v����B����ԉ��TܹuW*V��ؘ�+7o=Ҁ
Szz����ʐj���e�?���n���n0�����ꢴ�5JO7�Ì1^���Z����&<_Oo�i�J�vh�)}���~4
L/:�--MVE?DeE��~���C�Jp�;O�
X4�뽻Aj���cq�v;���'a�y�i�G�\fƹ�y[[�>48���ň�!q�����B����a��<1aus���2YT������_��,�t<E�����;T���>c<�|-��T#�����P̙?P!�lc�Q��5��Le�*t�`��Y?1���u�WIS$%ś�s�ʧ���U��1U��>�f���g�0Kh��Ҙe�~�o-����V���>s7m�c�l��Ze|�W��)I
�������ۺ,-���7#�@lU�F �Rl7(YST{Ęg7�?d���9���'W��OI܆D�
u����"�z��>Єs�,j`�JՓ	���ʝ;��CA�����F�L��C�C�� �'B=C0��Ҋ	5��5&]���	J�ڔ��U��ppp�RdT����,G�y�NLM.'��y߾u˪ W��C��_����A��w5�ME�
͂��m*�~�M���� ^�W�(q�z+ay��g����Ư��?v�y~��?��=0�`�
�/^�T7���J��s�������g� ]�z�W�A'��i��S�Y��t}�c�u�5V�����gtH�	�#�G�?'�	HI�W��/�#��*��"�����Qo�۷�˦�;gk�bDʉὢ�ן�LsS�<(/W|e�E�.��ZZڬ��C�s�)�a�BE+>��3����R_�<���1�X�!�L�-��0��cYX��Ӟ����PGc�ٵ�.my��g�|g֦�"6�*&&����'lnj	b��W����G��#��VOx3�Uh�
���1��#�95>L��+��9�����I1�ssKzz���TL�
�Dr5��`���Z��h�C�e�b�!��/|,�]�&|Y�FOgs���G�V�/o��m;"o��7�����q���N;|�.I[lL��4u��<G���g�?����S͔��N���¢�W��v��Hգr����󍣪�䎨��L}�.5Q�?�!S�	i�OMJ�~�w~�+KC�m�6mC��w�= 9�y�7��o����m���MC�6���5��>�p
3�ӆ��H���h4K�������M��\Qo�t!Z<��ĝ�:w5� ��p��[�5�Q��ߓSLRӋƂBӨ��)�?-## $(�p|��A�b�31VP`�|e�Ţ�"�3���;��4�(��bբ�		S27��_A�u�F�Hp��h*^ς |���׫1b�Stڀ��|���v�H�4R���my0Z��^��������!C��Z[��S��X���f�,��C��˔�7.�@����lx8��GdCr�����>0�/��1Y����>	����|�z{x���f��
�B�:���}ϸ�!uv���[ ���G����9-�B>2܊&_6�gt�!ƐvLhww�	�޽��������L� -��+{�4Q�[[�­<����8���Q~�������k�~|�c@({�70"��h_�����cc�u��`y��v��-�m Η.�� 7@���zR�'N�S����ukr�-Q�ܐ�Q��x������	�r��!��՝FNƁ@�j�����yX���o���	�뷬W�$6���f������a��s�pkVVU�`�����`c�}zQ�z��p�v�<�|S]{��!ټ%�:�.�!HIMR�n�ͬWO0I�UA�]Vr��r�$�����ژ<O�'1|`����a�5|�Lꡱi��˗G�T�_qWTD��f���a��  ִ������6&6�bh5�uf�4���*�vY������1X�uG{Qـ&c��|�-�WSTi$$%��c:y�����5��x�4��-^������x�W_�#X���l6M����ŋ�����%��%�-X�[]�܀[i�àu�<��q�kj��6^q�c���X6*:_}�U�K�q�	t\�ܹy�L'��wh�{LS������259{����r��E݀z��+��`#�\�D2UX6�締�猑�_M9x��Z�t��*RY��\L�=&&Yr6剿>o��J�zG��a��䴾�uR�ਕHVP�*!���Т�lc��*&c�0B�0���U-�?^,�3Jw8�L�ݱ���C�Bwh�q3�Avg�1D��WO�Ѵ-\�?>�L�Ԟ���2�蓈X4~L!RR�E����fB�(X����{�u��m��w�Іf��9��!KV>���^�U���4&�D�Z�*3	֧��Bҥ�!F2�Ee#�	D�C�%Jo�����WL+���+f
	Alޔk����l�^Pn�F�U/��_��8�ɻ���xo�]���go�y���F�a����5;�$�<�����֨# ?���}κ��X_��M�:B�O���E5pFP��EZ;Z͜ӊ���
"-�d�"cg)�ڷ������v�9��L���Ԯu)�y���֭&@D��g� �w�,���I=<6,'�:e��H���!cV��´���0��ڵ�VF�pt��L	��nZ�<'7�,���[��Z1�DH�X]]zr+�/pjIE�M���LqX�nh����z�n]���F��`�:=ynI��B�I> i,��L�mp: ��f�!^W�B�{�#����ޱ�(��a	�G�h;��>��׬��DK9�{
�tfnZ���-�U>�|Y��&3����+V�N�u��M����6U��z"�2s�H�jY�qDt�Q{��s3�i`dXr	0�A� ��<��lLۨ[&��o�ڹK_�Ÿ��zLk۰tJg��Oꆤ(LIOQ��uz���A�)մt��p��a�߼a����w�j`�s{Sq�M�r0�[��@�>�̈́��s����iCfG:�x��!4.S�O������c�uxT�4�6�g���9v-l����`�BN���.3n�JzY��G��n���R�>>~,��yUΔH��y6���QJ:��"u�v�N�[�u�>�%�
Nwl�&/�=�.z��ߓ7��E`ƪ��4ɑC��H�ae�L��(�Q|������y$|��0c^���#��}���I��ĩg$$"^:{���	��O��u��a�ғ��C#c�V��z�ݥ���gJ#04�6�*O]�VH�P��^PXda*Ƙܡ�g\�ujv��U�eZ7�^�=3��UQ�\�d�� � x���Th���
��#HV�l���Ҍ�����Ѩ|��v#�p�����P�E���ۂǿ��-1�!��u���^L��rJ'88|ai�CT�Y��:�-��[�-�����;\�jŉ	�u�m�7�f�c k)	U�̬����M6L�FF��]�1�}�0)vxg�nܲ�c�[sJJ���׾�		So�=#�}�WdJ7���F�j�U��Y����L2� I������/�yW�N)2�˴�̠`	Ro	/m`6�3́���&6���>�,g����̫m�[�}Vn}�R��ћsP	A�'DIvN�L�a�\hlT����A��-����F��	�v��ޱ�e����"��B����qB��u'&Ƽ¿�˿����S��g=V��˞�l޺M�6�Y5Nwkb���	jnTS 7n�K���ʼ�,?Q�施}B$$2V�*�<v��?|Hn]�D������~�Yu�}��\�H/-U�}�"(�%v�`p�c|�ئe��V�\`Q�N��GZ�ر�r��U�SER�D�S&|0����/��546���,%��\�_&���2;���W�RZ��ڲ�	������,�96e�(yIi�j�m
��G�ڢ�[��S��鐮�ǎ��?*K��6=�t]?n�3r��Y�ȑA�Qz�[[��l�ݶFP��2��
}T�.�>��
����lW�Ta.���//I8�����[- S�Hc�ضU6*�#WZ��i}��j�^NiL.hR��_�w5w��p�#��V��G���(��k�gd�_@���I�z���U�K�cYMdF�LL�Դ<�����eϠ'�BZ%<�K��[�j�����k�� Փ�����$/!iU ��"����z9�N�q�,'VO��3;7GB�C�a�On/-����t̕������$�i�P����J�Z��ΟW�.����'���0>wr�f��h~�'ޭ9zPZf?3� ��m��{�Eg��MS�Fm��1ိ��%^7��q������#o��i�������+����QoÉ���NC�inֈRhX�j���;�[	
�JSc�z���2�Q�B�4&�)�D�p�8B��k׮���$��!nۼ�
�f:\r���������ێ����_�gd|dЪE�3�Hefn�2��S����<Ã]}C���/4�xy?���`9��I���=��H=�M��m�1#݄'Dm7խD�qM�N�2OM:9k��ƦzK� \�vU�C���9�%�O$�����y/�kl:���g�Y��(�����m�2�b�Ғ�i]�"#�쏫p�qF�޾#�U���l�Rs�����d���n�X3*��㣒e�K�
LWg����U��w	�_�z�Qz<+��:�<�ёq�z`��s������Z��>�(m�]���%Z���������p̒˙�s_�r��`2����oL�
Lp-4�3��ﮠr� ;�K�?��&�||��v����Q�i�]��C#�E13��������{e��3H��{e��Ʌ~�Я�zx���?j�S���*�Ք����_%59E�*���4-�V[^�ﵦG�kVlc�ϑx�7N	�ƕ^Xvc"<�L�a���T5��$`�|#�C<��YHz��7�|�����~ʮ���`%=_��[Z�k=.>��c�C���`^'�x7D�-��4��8�`|R�{{,�����~����cq�+F�
\�fd!f�>��󈈓�0~�4Ͳ�h�{�T;������,�O|D���� n�R�Nxv����m�ڸIj�_������n3�q"�'����`uw�j�!��b�S(HT�=e���&9w�f�K���)�S�9TXV��(X^�ۀ ����a�Гr��}y��%Y�+�&a��(��ri�7�l�CF[�>U<iz� �,:_?��vǎ0NBH`��>@515�H;V�ɼ|���װ8�-��]S\FM���>�,�;-T��o����t��a��U�1��Qxd�3�O�&%�Q��6�~Z�VKL����2�Щ����`}]mm����j��<����L)�Y�0+����Q�Ya�ǰ�xz8��k$�3�����,d�W����s \����fB˹�
�۝�����6Y�G؆�� oS�H��
�͛���k@��Y �BC�ъ/����_~I��S���b��n���8���Y���%W����������Q����sX!Ϟ>%�N=-�����6��h�U]�?���iH5�g  4�",��Y�t�����8Q����C��o�X���Е�//+1��w&`���E��L��[oYk9��i��^���q���e��B�����,� ��|�uX�����8�����9<��N,Ӎ�����h!�i_Ô�����:|��y�l��{6�WRl��uYh�YS����޻V�hp���M��B	���Ojq,"�d2��<���A�;�_5���}h��6o�I_������s��=�?�c�ėU���,��>�鱸���d�ŗ��:p
��˲
YEU�?�[��n�t-��&�������#+B��q�c�z��u�����������`�rr��l<ͦ�ow�Y@�B���d4|��&ttK�-�������S����駟�������k{U+M9��z=��C��Ɛǉ�EƋ�sm̉F����la�^T��x�3�Q�����ܭ�cR7���ބ�0���2F]�
��\�����_��V����4�n�A=��?��K��t"L��J���p��o����F���f�]�5:t�l��b���[��o
"_�қ��9K�_/���Z�[
���������'G�WV�zxy0���a"&v�\�����,�sP>9���gsy������&R/����E(x@3�ã�Pˀm�� �����p��b� �i�`�8z�2���Et��$�|����PFВy�x�}�9(�3^v�t�:)t6cV�#��豓���i�س�U���R��l4�n?X�U����b�0W��ܞ��s�f�����2ߣ}�uĴs ����|#|h)�5`�!k�6b}�<�����m����ޏ���Y?֙{
�� ySD\�B����
)�F'%.6Z>>w^2�6ʮ��,�PZ� ���A�6I�SO��ד�fV����0F\oc�[U�965+/_����kRQδ�~IMI����o��hY׎� ��I6h�b�M-M��QϜL��֪ X�8��Pa����^�h�v�mD�z/��As~��[V��PWoj[�ZR�������~�sFG�L߈�m�7�811/���0y+�_���˯�ܡy�?'E��D�\|��7%.!��8�ϟ��}�`;8��#B�otB��yf
�4ʆ��n+����@�d<���ўh,w���wG�f?�я�3���/V!�G�8�\��X\X��Y�L0o��Ot� ::�����W_���,\�_#�Ju�$9>�H����<�

?���x��[ȁ��^����$).)��v��CG����E�!�u)���iq��eS̬�$� �@� (��L焹�1���zT�;Z��j�'���rN�:%���E+����ɚ,Ξ=+w�߳�FZ�^��vJv�	=n�� �L�S�=�͍������C�yIJ˰R9�iQ�X64���E=�7b�?������wX����N�o�a�n�C�����4�aM�S�\)�ɆI�
��}����~�����U�)"xn�B���4��������C�9k��q0�z� =�}��!��Ξ��P�)"�V���{�[�xA�.��_��˥�{D�cm��91��+��R���Zr�e�!�D*�C}]r��-���^���ͪ*�%J�L��6m庹�k-RJe$�1�p�QU�8���奦��`'�;-����$���L=������dsӇՔ���3ϮO�>&:V=��5w[M����̃��H��6��j
2�pմ�$R\Z!5�1i/���`��'/=�)ycQN��s{m�8!��r�$��ƧJ8�I6\}��m�|�3�yѸ�i6�#�����M�P!�	l�8����t>�3"(��F�;��v�o�\���6�͐��x4?�227�#������s��:�L��7$M����r���L���z؀.*^V=|��䔎`	���È+VV�<�b�X]P��l9q�)��Oh@��ol �l\����Q�l�y9��N������R��hL`q��U���f� �և���C���r�2������J�*�D��z������C�26JFj�X;;Z��;pPZ[�-�t���Z��1�3^u6���󌼆�a��Ǩ�J�1/�018��g@��Eg������;|��!@�d8��z-�"i'�ڇ 1� ���@#��˲��	6BF)�Y���7���{(�,�|�=���U�,,˷��-�Hߨ��!�z�A���-��SO����	�����L�drvA����xyyzy�>�{x����Y5Ii���30D������l}w��Q��(9�X�b�5=�?��F"%�Z������LϰM�� ���A���<\Y�,#��N�x�<�f.���Dh�����7��s�����g�VW��m1��ǃ�K����40�u����($"�ʜ¤4IK�ѳ]�i��]9�&Pu��këB%@1#�o�MZc�FF��}�J N�9�4�@�PrR]F�k�9G�s��L����1�p-�
6����{;����7��pb2�U,N�	_�Up�a|Ʒ��m�ټ�<̆�F�YT�������!��q��_},%�-2>�)��~��c���\�|2x���Z���l�}Yͥ�"}�EW{���w�7�`��#vbF��VXD��d�:,4�͸S��
�睪�.�����4���'��q�S0�B[���ޘeex�A����"��$&%H_�||����͵V116<��: �-����lݬ�*]�u�P�,*��$����i\��� ��1�JL��p���� ���V���H�&hV�k[��,8��3���}���ؔ.��322>�u�cc,���E:��	��ήu���#A�������;dX�%7��F���u>��s*���oY�\YYcP�TRe��ۚ�]*�����bnu�斖U:�H3�*eK��O�L��� �9!Y��'�7>1l�0M���z���)�=��=�;}b�!���"\�@��Z���T�;q┼��{��Ϝ9#;�_�<��)ή�[���PR�0%"���c'=��Y7 ���旬�L�\��҇�1�VQ^n�!���Q���Qՠ;bn��b�{�<�l�5S#r�r���N�ߒ�Q����'������&몆p���3�!���}�
πV�sm�A��mx�x�����ʊ�F�`����.�y��s��|�{�3�E�!F�&!�Vm���ha�n�%a
S?::nk}Y=���hy���!�sR[�&/��
�8��A�Y�V-8�d��㹤�pŝM�=�
 x*B��$E�P�c������bu�PG�)q
�@N��>ћ��F��)���n���h		>r��>U��R^Q*
l�q%����ܮg>wa��);����=(��6�)�\�L=��hF���b/b���S��23���	��l.עOrn~F=�����9\=���ԑ������O7!�m+�7�F;���T��3ʥK�LX�L�5������f��a$��ZyfRB0֗�c""��_~�+E���e+A�ڼ�3�4��>���cq1B=�6�@3�uu�m��h�?��?�؄dy������2��K�O������#�����%B;��l
U�Qͷ���֌��8`B��� U�q��&�g o3*t�~|Y^x���*���a4ά ���īB��*���ü���[-�����J�?$�~zI��_�Y

w���3�}V��&>�3�ʦa��"�I�?�/BLx��f���#��S���Z*7g�	��˷T[�Z75�����O%)%Q�W�b�f�~t��gٺe���G��e0���|L�l��F��5)����T^Z����K-�ES]u���������	zp�T;�h���!JhM�hFڴ������� V��;��D��s�I�|��S��k�3�T��Ĕdy�젣հ^��Uʕ�˙�^�=�I�Ь����ɠ
��hY�`��������Z��A��ʲǓ� ���F�V�{�seU5�E#�To��@�+r��=��
���M
DW����������F�8���O?�b�Ȃ�U�2��:�A2��ǃ5(9A�����ޅU��QQNC%��1���द����@pٝɌ�Vz�+���%�sr6Y��Q��i,-�Z�tI�����v�ٙ}�u�dJ�O����?:]�eL
&�RY`N^���6�-��$%2<ʮ��Y#]�>~>@uK��\��b��j��������G�,�i�f"p}�F߀ 3韜;'?�����~ �������o[��K_��:K���gyP^'��)�p�f�%h`���^&�^����׬xzz�h_�c��b����c�}��Z�/��r���Ŝ��f���KO �F%�1�D�8Uw��9v�j���t���܂�����7�96�}�N��E������6��
�8
�ֶO*�oL��$���LЬ ���O����6r��۲îC����i��g;��А	����a��N�K�]����ݳ�x?9|:���Wviy�15��V�7��6;�Im�|��G�@�~���0���A��(^��d�@L,
ain^Ν�@���c�Η_{U��ۯ��'�32�?d)�wUP�+������W�~*�ղl�Uk\Y�b
�6@(�j�a��z=+����Uoo#_/n��A�TTިM6�R�l%#+��$��-rN�륗ΨW�C*+�mzt�b�i!���"��_�v�kׯ�wץ�e�#���@�b�˦�>x`B�p�3��`q��sF=�`�|��ðq|!���E(a�(��iE�yG �oL�� f.x��e�Ŝ�� '�3Yen3&oR�yV7��l�a��D[O�"ǜ;�*�I�(��::6�fzn�;��dԤ`�3Dt��+4 ��(>�W�a�
�a��P�&&%�s���k���X�bIN=uZ��<�Z�M�L���G������KN�f�r�L.]�%s
��.�0��\^���԰9��V]^l�M���+#��ZU�i�p$�YN��/$�+�ث2��)	���M��,��g�[#@��p�j���G��m�pXx��%|�+�]���_>��kV��vw{Z�����{��u]g��W9thd�@b�b��%�0�d{my�;�g�{���7����ٲlI�D�")�")�"%0�	�@��C��ޜ��{_Uu7��-~`�޻��s���Ө�R΂�ʫ/�� v;�uB�6�C�V��S'��kX4
����v����p�.Z�T4E���;���z�a�����wI�:��f�F��4��c1���]��z��34��eS߃uj��-��-�Z��!��ݏZ��9��x��'Ō�8�[��]��+� �`��_�O~���ҕcl���{���x�����t/[K���XF�����/�+t���O�w~���d��*���j����N�	ߓ8g�X�'p� }�Z�|�a1�%\���c�q"�u�	��[L��Fd�	�W�E�t�O���Ƞ�ēh�n��ʑ��tjd�~���U�x0�4Đp�x�̳O�	@�j+�LG��x$Sɨl�"��TC���A�u����:�3�i�@��ρɂX,S0�A۠��DhK�6�F��2���(
�	߃�-%���BSI�\��Q^�~tʠ�|�h)ӿ����C=+"՟��k�&��� �p��p�"��3��3Y�����c�=��~�>���鳟�_��Whw|��Ͻ ��7�N_�◩���>B��������D�,�ڐ��ܖ^]�E�g,�sLBG��h+��c�ŞWB�j�	X�����ӿ��y�C>�5���[��e����6��D��4�iJE�0����I	���B�3l(�M,�����L(p�;���h���w:�N���ڏɦ�2_/1� �-Zj�bUؕ�*R�7y� T���x�U(�osH�̰���n? 2�*&E.��� l�^Kp�X�P�vz�C�f��C����#����]K��$�4j� ж�B�͎̚s�՚��.�%�����6�7
Ɲ;＝���/Ig4x���b�"�o��K���k_�����w�m��]J�lMjz�O�T���P�AE��2�-�S�����2CJ)3Q�5 �7]�`_�R�on��&�����#����^LP�P[aW��P܆� "���F�p�k�Q�`��FK܊�«�sl6Bb'' T�Z[!�puvj��P#�сF���%�������l&/�͖����� ���͵T�:�Mi���C���l;*F��=eC�s�7�	q���/�BJ�[C�L(��|>�(��p���9����Y�j�}�]��? ���vB����^��_}�����p ��+,X�t�F��,n�Mq7��ݜ�$t݌�Ø-���;��g,Ɠm�o$H�y~#4�H�?PR�/*�9���M��Q.�II�?��kT�-�=��J���Ǐ��ˆ�" ��B��]J�T�`�r<ż�U�WP��[��t!c�p�G.��:��[6+�,Ӷ6)����u�lZ�L9t������"\��0Q	kJD�g�2� M��+�u�#X����~��М(��&"\�Ӳr*�Fc��^hgh]�H�߃������VQH��+J��>�-cF��	^�-�c��}[
�PB��O}J���33�RA�!�=�����W~�:{�?�)m��f�.��Y,��u֨a��D\d :���9J2���)���~����Ll�6�D�`��5�+��!�M��wS�M���p1��;�3����(3B�s��)�-u���o�-�����1�S ��Hw�u��2���ݻ[6�� ����o��d�Yd�a2���A�4^�>Bi������^��W�l/\ @���0bSP�
�M�q�R�Xf�,]�D؎lZ�)��KA�[�4|ggWGT�<��W_��&	`)hjh,�O�87i@5��.^+��c����?y^�V�B��+_���i����Z�:��_xɕ��>��7@Ͼ��{��Ɵ��VбS�,f�xw��S�
D\;���D�et��`
�ֱb���h<G�k��2@��PON\T3©e�@�l��l��eͅ��u�2R7h�6�1)5+��7���Xx7���������kht���Lx^]�� �8�x-��l���M�KJf7
��:�H�-O�#4��'�؁Eh�`�h,`�><��`2��,'��0��Fc�"�-����7%AK���~��vim{���U���(���K/�ϞQʠѣ���M��L_���bmL���S/��*���\�@�K���t�bz���wz���e�e�I���
[�~�R����6�&t<-(1BX,1���g,� ��"��"���W\�Z ���̦pf|V�X$�T�h��㬹�1���֛���ECl2J�����#R��"ߑ���ɨ�
����V���?zJ(?��>Cw�y��\�r�sK~��'D�QG��bcx@Ƞ��i�\]�bvĝe��@LMN���j�~��[��fS> v*�eF�;Z�,+1Fgg�x��,ͯ~B��)|���H��� �q�e��"H �vP%�y�X>�@�,�`Rq���g$��|I�4?<��Mߏh�{[�o����oS�+O������>I��3|��X��w�N��{E���AC��PƢPМ�MfL��6�Jz^�P��r`A�9F�z�y�}fS��P�L�Kf�����M��/���h=�G�I��Cu����@i7M�v.14�#��׿�uY�x@�JryfZ�x��t
�{>~��AY� �D
�'@26^�%s]�d�b�=��%�����E�B��q�K���h8Tp �A��Ye*FN���>ѼР�^x�QI�Q)�'��ȸ�_�K�$oV� ������C��x�w��7ҧOi'� �aP�8H>� ��u}��/�W~�kTc<���y�~��41[�X�b��x���������SR"��%��[k��ݣ6Y�x�s��@*�Z�:�>�ܴ#�d>Б�C�Ń�'��H�$��7 �բŝ݋�?�݇�曮�A^����j�>�K�7��փ�U�H� ,C��~���i��s�3���xˍ��3::&�D�j��3	S��@�`�QxL4�)�$�hA|>�Η,],\�� �VD�!��1��6+�ா�JI����a�G�p9�*�l�H�����E��hU���^>���!�m���� �C�,Ϩ����?���I�ҿ�*��o�k�=��s�����NM����,R4Հ:��
1�]�՚�׉��Dr��I�I5�� W�v $D q;�`�}�2�O���X��PU�����=P���&�*��A����<��~��w�$�s֬́:n���� �i={j�����Ă{�O��OiͿ��;�]�~�$��Px��� ��^�Q����T3�B�o	��w�F\ s�^�6����L����[�L�PT^�}�C*F�6�a����%�瞳FJ���1)�4m�l~�=Ѳ8(2�S�]�@��$����%����0H�2z����g~B˖�����W����v��o��C��s/�w�K�X��Y֐��d �XJCI�����~�<�q�<G��N�tV��g�?��q��bY���h�<�J�@�%��ʖ%W�Q��0�5�����xL#��d�g1���y��	�O�G�\z9k�;'@��� ӏ)V�<�,�X,��O���+Ec�����顇�Ο�.�T&E �TAb���B����������0B	�|I�4j`�4E" �G@���i�jW�m;>��(�9l��N�V^h�x2)1C(RB�����RH�N^`�;�Rch�;?v���$�/�`��d�/_�n%|ƍ7�L|�W���on�������S2���n����̖�b�dn�1�$/�1�+�V�c���rϣ�kC�1�C��B��O+X�ua\g����ɞ#'U��יv�sf�h//�H��U$�@�H�YUi�Y����;d�prrVz���;N��v3{4�
��{[6�g��<v3�Z�o8� b���4c�we��⥔��g5�ᣏ��?"v����֛�K/�ӻ\KEx�g��":#�v"��ݩ|�2=�V6L(N-�P6���gdk���<2���6Z�t�R	���@�hh=o���<@۶���!���F1w(t�w-�����B��g�텃rk�<�oJ��<D�|�5z�G�R+�o�����>A� AO����|�Ƨ�8ݬr���d=���e���*��t�����k^��� ���S0��ǉ*ܻ��K�Wk��]%���C�#D������N�%�ڇ�����|��x��ϩ^�Y�#���b6E>U1��O'N�m��D70�B���wޥ�G��37)�'�nB6jlJ��ˬ�����[�#Qm�?��4%��{��Wh_��\�������C��R2iG3F������G�2K*�1������\:���&'��M����"X���eCAk�d<�^a���Yf��P&s����9�����<^~�Uz��'�K|����
��}�6\z���?��+T�Ts3�e���3���`"�-$<@�:y�
�;��QC@�qڬ��B��	�GDb�nNͻ��&�-�'��$�e�ԋ^k0X��e���袂# q���V��5b6�_�I�sz����q��^��ֻ��K��h��ߠc�Q�����B͔�Q��p? �b��?/9HG:!��#���_|)���
6}�3
���~����)thr��}�_����3D����a�c�B����F.L<������Lq0oP�Y�s�l�:I>���n�2�\�`X�<�������#�B�\'}����ٝ������o}�z(�1@U�-��s��7X����5tMGm�?Qƅ����{)���9�_^�R�XRw�!�gp)x�Q'����C���@��v��7��/Ȥ�Tf����h*=t�=��c�λ[���u�'���(5�_yUZ׻:r�b�R(��u$D�t4ZJ�B�"@�d8��H��G��t0�NG�d�!4��ڹ��瀍 ���@ٸ����T���Qq $�rB(^��� �c�R�����+�0��u�8����w� ���lƑ�A4��Ra�>~��|�u���'M$�����O~�6\|9��Gz�����tr�@]}�¤ɩac�y��*H{D$�*�vec�O7 +��M������+���^Ε^��*�*P�+poF�тߨV\�z��Z���	����]�h��zy��8L#c��4y�Gh��}�}/]v�G�^���r9�_��~�tx�)�aO*�*�L����.$����)�+ԿLm�AL�H*&��**
7��=;5vg��0x/>�Ρ�C@�����D��1�.{�C������e��HǻAH�wLŐ�
��d��M�����}�����>J��e�x5�ɟ�g:w������c����ǉ��:bv@|OƀMu>��TJ��O, 	(�'(6 ښqq�XҼ����`����؈g).���+��~Ih�DT
��-��I9	��*�t�Pc]��k2�Q���ʬOQ�Qe`?26K�S�`RN��A�׭f�t�4����k�clF121��	_*.5��(�_�P�T�QZ��?����5�ꍪ칲#���������Ih��C��%��e�O�e�P�CAB��	3�i�:ILh�V�>W�7�p��i��$?�Z
l����qߵs�$�����-7�&c�^{w=������LF�k�r�K��X������ 0숴��?l	'�
V��k}�H@�����:��i{�`	ǘ����A*�Zj�uZ���&�|si��:�d�_�rT]vd�R
hɲ�TgM���	b�kbw�Ta�<G�cǏH���k��}�}�_��W^�=���I.B�B�dP��� �7���X�o+��3ԏr�G�)d�)eԳ�x�&��8��M�vH̦97zO	���S*d�{tߠ����K.dsw�t��1����$�b����W虧"��-_E�������'s]�����η��E[������cA�b���.���*_�
,A�j�j�mZM��n�N���������Q~::�ԐN�H�+��b1>�����R�@��'zdO����x���bZ��_L��X����emƞb���5*��X99IçjtΊAb ���]�g�A:w�*��+����ϥ[�Y�i1�!!��悳`Yq�i#��0j�:/x	�}`�|~@�:Y�C�E`��[�,�UwbR�/�t6�Ӆ鶺v��`>{�z%���%L�В%�Q v�3R`��m�z���->@ř��R����}��+h٪�h{�O?����kt��5�B���S�-C2�I�"�Kܡ��v�Z�P���Q=1����w��u����\mj��>tjg� ��M{im-x�@��D��߁�H�@��h]�G��`�j�8!��z�jr�2�Z��z:��/��{`�q@�����S�3Oe8a�I0��������xW�֮^EKhl�*M�>���������=1oh���λB��'0��^`�)�=}]l�V�P�Vq��ӊmn����|��aJi4p�i(�7���4ojY~m�Q�>�\t��8�<��!�x�1��6�#�	�àiׯ�@��::������o~�Qz�'?�]�OR��=���Sy�ݜ�O�5�OIO�	]�|L%���r����F�4�3��bi�[���H�o�6ޠ8sl� 8�`�b����2 S/*�q��8��v\2&Z�|��8��4���\y�Ŵv��`	�ȥ�����
��ŗ��-[�go.�'�e�U`-��wov����j���3�齝�w�qZ�x-�.X%\U�����cP�!���������ݾMZ�+0�$�BS,�Tv,�<=�]�:,K(gy�q���v�x���P�*�51
�c �_�j�$�����$ݐ'O���M�+1<h8��ӟy��`-�t�8��O�ˏ=G＿���9�p!Iپe|ST��Mcĉ�g�y��Ii}l��rM��]C��l�w�#�H�8&�@N�i�3@r�̦0�r}�u|��-.���a3�m5�,���r���n�/cTh`ȧc�#��s?�����A��4�ul���i3��ƻTb��X�Έ���-ÛT)�gW����Ȁ%4I����l�ƞ�fڰ~5؅RD7�n�?~�A�^/ZD�֞+4���wn�139%�B�D��9^!P`Z�Y��B4ա���$L�0�T3�]{���dd�̘>��P"�9N�w�w�&ݣ��^#<��|�����hh�@���N�O7>I�����}���G��x'�Ѧ�׏u�lpT��1�:��؀j(��LI��m�pA���l��V�eM�z�V�yF���:��b���AVS͉>�
J7���5z�<����*��ӷ��u�~�n���i)Wk|�b�n@���ㅫ���\dcb�dV0��
k�����˚odz�&���6m�!�tW_y]�ћ�a����x���k�B��#Χ�\|���EC��b�q|6# �(�`��Ŀ=�́�u�SV�dZ��HG���[��jh�+����9Fp�!�(�Z��ֱy�������l�M���M[���쒉��� gz %�2 \ORZ	W=V	
{q�E�ڵ�"�?-d�4@���&���j40Y�
�ڡUc)�:k�/L�ި�l
#��M���Uh�e�d��2�����K�l�o"���+�c'�Le� X#�b@Ϙ��I>�Z��X���6��E ���_���J�i��5��_&c�ff���#����lv\���@�_r1�bp�I%%O�h��ol��t&p`�{�0h��!o��)�>@42���)�J>)�NJ+>4^��I�j-�Y	
_{�e
�Y���c5>1Eon�C���� q��3��9Jt/%��}�sT�1����P~ႂq���H�\#P�tlQ��<��}l�v�j�B��hᇡ�3�� ��
�K\a�%�*H��>�Gh��FR�3@O�-T�L��t�`�/��_/��1k�	6i ��	��P��Y��@���3��#�5%x�p�cp,�4Q(S.�E]�>	xb����=���s/n@���fՊ�t������/�PH\����f�hxd�=��7���Zq��Fr�ֳ2�%!I�����'�	�I�!9��=�&n�/?�i�l~��$����k0#(In��=d~=p֑
c���2�'�
B
V� �hT����.#[kb��,��(V���0�m����J�εШi*��F2��Eu/�,�)��K��E�B�jo� N��h�ň�Z� �<�HLWA,�ل�Z��%��������&M�!�Q��s�`Ap�����{��*�	X<�E3%-�Ma�4�\��!���mC��m;��S?yA��(�Y<�K�Y���%�[���>"'�d���xC�7�Q2|�oW=E��Iw6"
�@8�g�:p�(��O���s�g)ɂ�Qm�x7�/�j�J�'���Ћ((��!e������m�тƲ��,�2�5�$s�5��	�e��0U�V/�1��9�wX��{�M���+�8�#(c2Eݮ���M:Յ�)whU��ř�o KOLL\Lrth�b)�5��'���}!ocE~sa� w7�JUGpNx2�LbL�H6OB�L��t/oU�vY��&͜��K42y��Q�2	�@A���� =�����9T1=�$�H"�HyQ��P�R��(��)�� (�{����9�D�m:)�k�CF�ŜH�hPו�����VC��,�
"o.�b�V��;tf���lTc�"����z�RZ�(����z����sc����HWD�)�ы�+�1C�
�aC]��ɍ;j�bV)M+
���@x㮆(�g]�*�sI1�Y�@�]����$=��#!�@LR�� :��X��ޗ�B�d��M���e�M"M������:��&��� �[]������S?�3@>4˙�a(��>�H_(�R��y(MX#�6�@����mf-��i�{�Զ-�KQ��	V�i��c�E�,G�c��Vk(�O<J�L���Qzd�qq��6����@����
Q6��:T��U��:�0�A�Az]s"셶Erm.�����Fo��XF��X7�PV2(C$���O���H�'���2���Gk�*l�3r ��4�����6�q�9GA��%P������S0?��s����9�l��7���}���H��(ᨖm]/��9�����" ��Mm5�w4?7}���k��:0n�D?
���	Z�`ч���.X1?P��]d�t�j�9���� l�l� &B������.r�~T5�FR�ࠍ̋���C�9�<@ng/\�N6�U)Q��dxg[��\]VA0��V��
�C���7:�ZB]�-1����O�u���Q{T`-Zkpt�؏R'4�Vտh��=Z+=$m�4CS�E!�=-�)!�OP���h��8go��p'�;|zS�y1\�/�g�$3�MM��m��\>��1�VO�U�ZAakV��Hf����zU�9�˅		�"a�bosQ_'�O�RP��I~>���N!m�3�p�sk��-K'C�p:Q7��wC�/�j�B1Q�����x��R�PȬi�l�>ڴh��6�b��vϭ6��XH��c��j�-�{����k9��y��]���O���zz�J!,`C6�T4F��so"�@���dOm{Sk�F�*ڄ*l9q�9<���Uv���)�Y~�'��<-b���W�W��I��>�p�'?a�D��?!4 ��#ω�t���&�تn�z]csB]'*r4p��p��1i�$:F��/bq�������&�����4U
��{¶���|n8/�M
d�Qўo��Q��QK!�c;�b��4�F�����LIa�<�@���t���.�s��pN�;+\1c"B��$:�������_+Rif��)�z�Y�c������<�^�\�><���t��1��i�f-��t�MNI�H��8B	��hژ��&��rԒ��i��d¦�R�����y!��r���9�v��)�w�N�- ^�,�9s�N֦�;#�!�;x����KZ�����迖\�fUX\��5�i-�T�8fꡬ�ͪi qިDuX{u�y%�FeZ�Y�{��O+;st�G��Sc���KoR��X��4�ڂoBW�}&�`�sM��:W�6�#��f�.~x�� t\c�5(ڲ��i_�
nSE9Z�+	���m�rG��i!�)i��8�s�&�E=�&���Y�3�9��5���/�?�`���͟�@\èvj�R{
�
�0������i,��gj�����0"�h�n65�T���~��ˣ�Q_h$SID�{��?B���e������s�^����ݒ
�\�ݫ&J6��1�m����Kh�_��>#������m>Zq���[ׯ���7Z��������<<s�}.hoj�0�iF�U}�t�K�zZ��:����`�%~�/ ��m��N�<!k�{��k��asK��՗�ِ����$���.�V��#�S��ɟ�&V�6�iO���G��:���*&6�q���^���s���>J9���3�3#/Rs�ڵd��ܖ�W	���RQ����h�Ē����y��B�{�XX�MPs�Wk!��w2�l��皾���4����z=�+�OǊ'�7�V@�N3���`����p�Z����q��	X	U��.��FM��W]'��|Gtbx�܌���ӆ�����)��	Z�}^b:dx<�D	O�@�wgLlTK�@u�9��x��S�����m��Ń��B�M�Õ,뭪BQЏu5ެ�~<b溭p5���$|�f�[�371g_��{�W�^A���B�2�ªV/K�ᶜ��mo��ʌ�!�J%)/I��Ck6\B�׬���S���LwyD�ӛo�+e� ͨ���l.�W�p�K�#%jC��6�k<H��׿;f#�S��J�L����u��v�x�=4�������D�Ɔ�Uq[LU�M*z?&�᚜kH2ĉ5��Gp3���Z����{c�$��D/+���
��4SJ��h-�o��ӛ�d����-ƴ�`E6�)� s��B�غ����߁&T=�.��>�?:B;�����q!	H�����MO>�S��8._I�l������aҰH����Z�F��\[KW��h�+��P=KI��?����ɵ�.�hИ��̀��������������.\)K�k�P�N�h�y[p`\S�e)��vDV��I�ޭ\�Y7�����ؙ1��2-�b��y�*\�V[Vw�G��8?l
n�Y�_�3�[��'?��R�D�>�Sںs�w�Z!��w��ڳ����z����b�Ɏ$vØpl6X%�u��F���X���U�sX�s#\��w�Ѓ�/n~��6�2�KB����hdH���j&���x��$)v�Q\h7Z>�k�p[-a�و���s��N���� �Ms+0�Vo;d�0}�^�O��ɖ�g��/[DB�H��h��������Ys��
U��E��u1������x2���A��E�Α�,x�,@j����+�RT�T��t� fC-����uv�<jb�V�z��=X.0�:������-I��B3k�/~Ska,r&%�/�����c U3Y�fC�uFĬ�9g�`��h��&��*&��C6��b1�D��XC;��.f|~8&�����x�V==xOWs��5����8�ltR$|���6W�E�9�%d�9��N���4�%���'�)X+���S�[��)�$��i���{I��J�$��'24fBpZ�Æ.�uV<�R�Dh�ɷ�L4H#j,i���#���JU)}o�U'�4;Es,ضo]�֘�{��#��u�>���-��QO+ҙ]��V��\o\#�q�c
˃��i�C9�h$N/X�t�l���E%(P$=���3?Z�-g�Y���0���S3i��w�J�g6��fLdfb	�����:裺R��д�i��+0���.iC�Y(ႆ��R��j�@�
��j�b��'�^��C'4T"fds�"?�aS�����`XA*�$;�ıB6�@�h)k���(�g,�/���`5��@jV��,.P�Ύ����&�覻�3T�d*XZ�~~�tU�F�vz��w�(���@]���Fm;��RB�5�(���k����>\g�?6�26���k�vL�@p�Q�Rd,|X�*5�&��8E3I�V���$��6&D�TS' �0�-�!���S	�g��#����s��\.O~�L����)!�ŀ�reJ�0b�u5.�Sꮤ� �Z���\&���D3�i��9��Ñ��IÈZ"ֶ�<���5��E=}VPb-pCㄾxrв(_��8C-� ��W��5!��~L=����h2Τk�30��d�'rDm�R�#�
�j�zz��/�qt	�b5�x6,w
��ހ�Np�4U뉳3Ws����p����ba]����%C���e�c�}]����,XU�e��>�8���WOOLR^:�C���{���F��2�eS4;r\��vK�F�� /^�l�ě���'P-���>ũ	�9+|�y���嚪A�����DJ�M��X�ԯ Qp���V�4�9r��9��M�l� 0�[�bc����c�!k(�� �-j0��>S��FǙg�ک"k�� �7xm�֦���`��67Gx�z>��{O'�ss?�>75=&�Y=�G�)O�����'G�������/����'��-�Ks�4SP��O��?g�39z���7z\����0u���s�Mt�5WS��bZ�l1�0&z����M���C'���gV��b�l�X�Ăg8��ϯ]��n���󶛵��Ҡ'�x��y�9�(�ױ��h1B�qrֳ��V\e�墷[z�P��F�%r�`(<U��tZY^��Gy5)�ĵB嶘�|��X�m���:�	GN[���*X��3>�vv�t��0��y��¬C����ZHI[af�:�)���:�̥x�ج&b4[)P��k��*��x��)vx��R�r,t���_�;��Q71��q�L���n������7���c3�� ƀ*��5v0\ntB���c�g��`�V�����͎��O_~�f�c�L�y�i�dR�|�o�g��ߋ~jI�+��umD��:���`B��)pUqd��q��M\|�\W�`-��N����۠}�?�`ѡC�D�%M���F�O���t��w�t�B������& �r��6	��P�qgQ�56z��ѕ�_D�=��!�W����brk�i��u��a/�V�|>CW]v�u��Ԩ���������?�t�H�V���}�W��s��o|����):15+�6��Xg�7[lPcz�v�)���^>v�~���izj���?����~򋟧���B�d'_C�pC4�AJ`,�M)[E���4���4_�"��{�Z�⹮��m �!��k:Ѿ���sea>یh���!�z3�M8�܅g�]�kN�8�{]e�s�����G\�K��0�m[ާ[n��M�-�����Zf�Wa��}Ǉt�%�	/���/�d=��Y�ds������}���	������c�8]�����^��FEkIZ�X�;K�C���u
�K�����m�K��B�'gg(�ꖆ�f^�9Ip��,-<'
O�R�ì���B~v��]R_ґ�M�92�
=2O�����h�w�kj�ӂ8���n�)����������d�&�%ο��a��@�Cg��a��_��k��B%��S��u*���S'Ghld�ְ�������^��+��c4ujZ�xeE� �ӆױ���[�b��c3���RU�_=>B���s��� �,yZ�<�̔��,ߑe��K�z ��5���߇�:�7{�i��-]8�L�6�(R�l�y��*�#+(u���w�n[�C��Z��v^A�b���06|cr!p1O�"蔒�3@bn�8����3��+��F�?Q����a�iZ�+���5sź�$Dg�j ��e#Lz,haM<&;�<�l���g%]|�E���Mt�eW˼�����ĽɔP7��V���w��)�f�C�3�S��Q-�*��J�H�4�ש��^�2�$}���Ӡbէ��QZs�
���OP��ГO=-����׬,�8��tט'q-�j���ޡ�ٌ�B�r�U�����k�����ؼ�P0y����f�W��4b��u(� ����9��s�)Wy�����h�v�D-�AK��
Ck��"�;�s-,<��([_��;,�cP�����R9���p���[t�mw	����_�k��J��ko�A��N*UX�ju! ��
b�$�0�/���_�W�$����<3��.N�t'eso<An##%G�F��k��E����7	e��қ�i�ֈ=�Wi�HPl&By�5� RaK���\�^x)���SCն�(�����#U�a��j#�i���X!2�~��4\mn��gE��9�i�Ӏ𹏅��\�9[��Wџ��oY|�L�øaNVCxLQ�f�j\�K�ןG��Y:6|���2��#D�Ha�G��B����r):��\�ԐH9�]ݒ�9~�����޿�����(Ş'�w��=��OC���#G�)#]��{���4�q�{~�A�m��v���キ�f�u3*�ɵ��,���JƠ�ֳ�o
hL��^�hz�c>xg�q.Xl�j���Z=2K�t�c�xVk����ل
�O��d �dNrqU/c,l�jM��Tm��h͚Ut睷J���g����]<0�1p�=��G[?�M�_{�x����OQ��wh�*�Ӵr�b:w�j�^!��s�2�n>�I���X2��Y�Xa���q��������ߗ����`���y�P:�fp�hYU�4�4j�M�u]V0袲�9s������M03��4�'�q�dUG�Yd�_ۼӱ ���D�m���Zk"���)�$�n�B�`g�ӝ��G tDȹ!�T*ϰ�I�u�8B�332�TH�ٻ��߰����~ؾs���t�`Zh�9.�7�~�.��J��o����6M��5K������&n���,����|!���kJ�7�-��;Bg�ۓ�?��ߧk����~N����Re�T:�\��/'�_x�%^4���z��M�|/r!h6�%�1�Ӳfa��e��]Ȭ�g+�[��r͆	���7,t�����?�5�g��Z��q�@�}�f׸��c3Vcͣ�Jt ���D?e#}��O��)Vh�P�͑[���)k�*l �;����>{����˯����RL+pbV�"��wh���B���&x�lJg����}�.X���3�t�5W��\�涃≜ԙ���}�^|w�Bl��svҒv8�B���K{��i�V�+`^��ȕ�?����?p�ɤv�&G� լ��c>�R:�6{�J�1��`Q8O ZU����羧�;Z�7h��J���>Ֆ�2ǅ�!�bO��Fr)�22*�B������?��&&��:d��]�@��r�ƾ��th�A����К�k)��h߂D������[�Q"7@�����N���D��1X'o�r�>��������N�	V�N��@����N���Ƃx���]�V�aٶ*�5%�g�o��y���>�_5�S�b oݶ7-d
zk�tt]�x&����W�6#�����)��4S�-�`ӕ�wH��'�R*��r�H����ѷ��;�=�<���X���?�*`�<�?߽X���������9��MH��ė���{[鵷�f�hP�A�7���A���;虗^��Z�T��5��VXk��c4S���}�Q���X�e.���	��Y��ML)��"2ڪy�6%s&�X��F�O�E�m��)d*�9:f�C-�i�8+t�a'S6�h$�,��3�B�̧J��+�0� ����`�ߔ!=�F�-��]c�C�mY	�w\�߶PsL^�����lZtI�
�B��R��iU�r�dC�S.e�i��ץK6N����<��Ta�����)%�`E6� �-Uz�ӯ<�YZ�v-���HϾ�s��֡≸K]=2� ���K�5UX�Bf;�V��+�G��ǂ���J�#��}
Ȗ�$b����jy�,m�˵e ��4�Y1�h�	�xU�!ē��Z�̦3���,�0��B<Q5����^�i�����B��8�hv��(�M� �=�u@62�\%~����hF˘M=,�S�v�h��&h}��oA �x)�AJ��x��{��� �*C���ע���s���|��l%�I�n*&f�%y3��C2ɢR��3/l�%+Υ�����>�ҫߠR�Dq^#tl7�x:�Ԓ+א .B�\�/�`�V�C����aK�A!d,pl���	����|�*$M�U���qYoOL��c�ʳ� 0pj�q)Rb	��WA����ar�@@���8B��V�x�~fS�S�l��KM4�lh�R�H�j�CvaT�i�dǉx�����t_����Jhs A��&l%v��8�ś+�Ԫ�Z�I�$Ϧ$�YX�)P��xQ퐁�P[�u��Ed���ǿa��.��@�|G7�����?�?��7yS?�y=�r�c^BJ|3٤��&���C�w8qdn5`�j����>T�Z��j!k�5���A����f;��oH 9�L��j�D��6p�"9�M�Ϊ^m+4Q"�NX(�x�/f�Q�!���C}6�Վmdp�u{�@�>�Q�+�|O�B��Q�@��Y� ���ʅ7UF�A5��T&#5Ldl���1}�Xװ�o#Za�\�(�6�Gj�K�^�(�c�^�_II���|�I�2��Ԍ�3`ҫ$�;�3d\.�<�R��#�U1G&��q�{��в��;<װ����9J�P�Y�#q&\��
��N�H�M�@�L�/�ɣƶΐ@�L��~H����0,ȧ��#N��uvW2V��R';5����YrMձ��!/���}��^&�dh~���<�K�k8����6����$��ӌ��4��>K2Q*�?�w�*jÑ�l��dc��8
z�ۢ��!vj��[�IF�8M��Mϵ���	e#��lrrf*����9�L`l���K�B��9(��C��R��v��H/b`ۯHcEdU��A'����m���35	N�m���ݼ�P&�0�K����Y"�1�@�l�'��5�b�^PڣN>(Hke��J];�j���?�ae��'�a��ę�a���b3Y|G3�iV�H�V1�/$��1|��_.3�@p�D�JIf�)�m\N.Ʊ��s^P/��,��@
�j����E@�3^م��S�,9ԍ��F+T*d�Vf��<��EF���V{u����D!��L[}(�<!Pr?�]�I�,�"C�`��C0p �Zy�#ѓ�4y8
[ۻs��	B��n���R���s�����*\�T�h�܆�]<�&1G�C�OY>l���q��R��cy��:)��&P�g�=��]J��Ar��0��pc�����$�g�����EB��&�ǟ�F� �F=7��um�ʲ�/�[̦#!����t�`@���%��Р�
4hU����Ϩ�߶9�ބ�Iq�XVB#R�L�0�Ykޛ��v5���I�뢒�m�B	I��<���	tؤ[�R�q#(�-�
�4���ze�	l:F���6��ֹ^30��C�p�P�C����@k����t��c������:M����QJ��|�"��[E�])�ݩ�	�����]�%�֙x�Kg�$�`9/ҏ��h�%��bU�T��/�0���k�'����5oԊ�fo�K.��.�������2�����ct��0��}�������k�|��I��|:�a�o���:���  5�IDAT�k�e�<N��\�1&�H&2':!p���5	��e�	M��1��k�q&�VB���;�{A��B=L����J�����Zi65��(�Fk��mƑ�w��Hd��>�
ikWh����/J��ʳV���R�4A��l*�t�W�}��M_r�̼��YFo�`�]^�C����?���cz�w��g9��C�{�9D� `��\1X���j,!1��UJ�gPg��ڕOSw6Cc#'��t�%�ݷ�B=]2�avjR�.�@�Xᓻz�-]<H��/������Ghrf��_�Un^d�U����W�q�CN��W͇�������-�VO��73��u��B�θu�<�Y�*���I0)&�v�$�	BS�ь�|R4[`}���TJ�ݖX�c;��a4��Kٟơ�y��Qu�&�u�e��ϲPud��(OҩchŢ~����7]'�15v�
�޷";XS#$��7��O�{]q�%��3/Ѓ��*��1J�%x��T���݌�1�g,�s��,�W��6�#�[+��P x�u��5W]B��;�Z���R�p���bZ�4`:���\ͥ���E�x��"�Q�^�.W�6�̢��z���'�&Q�6@iDfq%L!J�+�����F��aKC�@�O��:�Ơ��1� ߋi�6��8[�/�I�@�{�(;��7��VrZ�i��j�U�k�ϣZ+�1�Ѓj(S����hҖ'�:�"��@����-�h��љ��n�h��!Z:�M��o}�.�xՋ�4Ç_���>keG�.�Pf�
����}���~�kP'c�o?�(�=r���:���(��V�Ĉ�$K�B[��<���=_İ8�
�b��u�`���\��ןGW_~t��k(���a #:se�|�(h�g�����^����[���7�F�2k�4�ϘN(�#Nx7�j	j�b[ m �@�t�	����5�n6W����i��R&Q|^@�JY�IO*s��w.1:>�?"�Ё�!GCit�0��`�)������r�B�a��'߼��<��8TL;�a��$�$#i0&^c�zM*>C��f����z�b��'>F�[I�G���%0
�4�Qu� q�o�Y��da�Q��C_��=r���Ϗ0�9B��&�%e;�T�<�+���1G��ǆ��E�AШPw>+C�מ�Tkh<@�A��c�Mc�,GP���[ɂ���th�|:qd?m�u���J�bґ�ש�fz��`"m�P�x6�������9lr]rh��&�9Z������I�n`i��5�^�VԴٮ_��ɾv<KT���0i��Åߗe捲7��	[ Y��|�2(���a��H�#�p�̰
~�������)ȥ�T�'ׯ�m7^K7\{%%����Zw��e�E(]�[��.��#?u�mt��1z���� ��Ĩ�Zc�u�o }rf��o�u���d3	��$���������ES�X���&pb�hCk#������j�N����5���Kh��8���/�%��:�v#m��M�û뵊�,���З�Hb7�E��p�r��+����G�Ml8�!�x����� 8�@ӆ�aD�j����t�4d�J:�P@�b�1�P�Z�&	���QD���q�W�1������޸#��EGZ
��Pz�F]&5錄I�*Aٔ#����h=�����Y�<�|�1��S��iF���AmPA���T%�^C�v_�ґ��i��s�6�2/�b#8y�������g��g�X]BP<G��$�٣�g��%�e8v�0&�ñ��U�iO�I���Ǥ�AǗ��]�X2H+W.��#{x���S2�8��:#&4 �1t��LROf���{:|	9���A�0���S�j�GT�i�2B^�t:.Q���tT!T�D�������13��)m��" 
�>dٔs
��&�S@ z��K2����$Y��Ų�%L+�?���H�U�*40���'f�H�brP�(ܠ|�(0�#P��/ѕ�������C���l��+fLK�N�@�����g�.u��ʣ(a�K/:�n��*�y�u��*U��vW(D�r=g,|�-��!'�O{}=,����IV�劘.9G��0$�D�7�D�e�;g�,�|Jװ����>��w
qr�(s�(���au���d�����)�U
�_r�T/�x1�,����$3�ꗪU�/O`�㞉��)��׸hE�I�HQ��\ma�Ch�����4_Ogg�Ҭ�fI\
�)�3z�;idb��$�'� #0���V�X-���,)�X/JS���C�;�q��o������CR\&�ńg� ��Zxb�~�9��B!�=!I�ȁIɬHm�RGZTH�`vk�\sB�M�Y�5kVP������`�eBY�e�{fS�����d�Ɓ���g��<����� ����+M�[��~���|�����#3|3%���Ӊ+�Ib�����
���,�� �O(W2,2p��$L~^B�"�<���d���ŋ:y� -[���;�4[�H����2$s%S�h�L`�L`�����5:9"]�ld�O�=�k��q�J�Hu�őb7���8d���ϫaZ+���)�f�ba�ǫ'�������3�|
��2�:%��pH<	�_�b��@�N�E ��y��*^x�1)�7��<_��M�4���С��5hӠ\��CaB�2�0�9K������F�I�͠vӌ�j2�����H�x�5�v�2�)+�`h��ʤ�S� #���ϔ��*&��ڶ��w#����3,P��a�ki���ɉ-죎������O��x���}�92"�y(��Iu��d����i���t�9�dP8Xc��=@GO��_bӔ�ɩ�g��MVxA|��S.�fYS��e����z��!Z�t��c�!���_�Yh?��iI6''�5)M��k�ko���[�������]���C?N�������B�. ړ n�)O�80؛n��,;]%�>8�	�·�E�U�qUCJk*��,-y�sb�x���t�����˳�vj����!c����L!�b?�����Xx �|�=�YZ��)Eucc���U9q3/�!&YH���L��τ2)Z�OP+���MG��b�B#�Z0�a�}Oƕ� �a/-��e}�R�șhQ� ^�j�q��id�"��V2��b�*u`]��l2fƎ��(�`�5M����d���������Wߣ����� xeV��OT���4����1���~���z�MD�:Z���75;z�v<�� ,��zMbPY~ry.�K�8N��m8o-]z� o {\c�����=_��n������6���.~����}`:j��5l;>�1F�a��H��.��5?0�PL�T�k��p?4$ Af,�d"M4a��bh>�\4����ET������txF�����bCj�E@�Um~]&�g.X+C�Q ����BY��b�x^�?��"�S3Xō�h£�=6&8!f*!�#�&�'����º���":�{���
5Z�l?7K�V.�����i����Ok=�I,,�.,6]��8u�^��3���H���c��;D�l8��{y� ּpɸk*6]��#�T���^6q	�Ѱ)�b5;1L�ޛa��fS�A˗�(�Fc!�y1����Y��G(��!�������$�?˛���ї>�E�ؽ���\C[v��S'�kp�T#�(U0�}������/�R�&'�i�P�ZRoړ4T��R���%a�)!p���*8ChQ�295�V��8��bV��NP;K�]�ر$[��8�L�zww���O���QqQ�W2�tN�(f#˨S��'�,u$-��i*1P�e��)R�Kb@Џ5%�>�ʱW�S%�;�W��8��R��r��V1^�3�}�7{u��"T8���O3,�1xAlZ�G�l���"ԑ��#��-[���%K�q�?|����&h@�?�a�,8��v=�&����<k���=t����`�������ALJ07����׎Ӳ%}��5�у{��j�9�ݰN����4<2F+�]J�]|>��i��Ka(Dr��	g~M�/._7X��Y��w��:�bM991F%^�T��.�W�'���奲��^���3�7ĥa�@�<9Ja%�	� '�֨{��v� )����T9b��!4x����8�޵��Y��O�$����?`��������I�����f:�XmС�'� n�\^�zE�����WM��s��R,0f���W,q�����N��=�}��}Z~k�Dw��lRf� L�J2I©p�9+��M���	���a�]���yz����g��}{v���s���?F�w�-��,������n�Z��M���T)�i��!���kyNһ�oea�fݖc-��S#��xd�x�rlV+�3�g�޺tު�2f;v�k��x���a�z����|].��6|d=��[|9Jgsb����V�T��|T�3��M���N���1�B̞%�8
( �j���?�ֆ%$����:�|��R|�����fK�(���"�%�b��g,7�,�TS��3�.�S^s�t�"u�d8��rN�+�=�&<�e����qZ�O;w�0e@�%�M��.hHes3��A�#u)�M"pY��ﲐ�VI���bqX�O�4��i���S�I��	��!Ց�MӚ���8�4q�x�'��cAYGs��0�4�}ϭ�t�Q:Ƈ��0{���dc@�r�v(����Eڳk']s���=uJ����u�f)��b;h�Q<x�H�3 �%�����c�O�	��_����IvZ�l�C9�Z���P�� �#a���l�J��=v|�^y�u�����t������9u�N��@���h<�<6����#�������{��~�}��f�G���6�^�>���*F�B[Z`R(Rx�DA��_ڠ�'O�}@w�vK�'��8p8��F,`�eȅ��g��ɧ`�ì�={�I��N�|)���p}�#�&��1Ʃ1�j`�/p__/�x㍴|�R�`A�[s������y�RbR=���/�R6�kl�=����iժUt��Q:uj�M2z�������ჼQ�5i,ߓ�8���S/���I��CZw��b�
�Ŕ�5:p��~}EO��J�V�	>��uhd�k��B��a�b��FJ�<���i�p0���Θ�ZZ��@2���J Zm�5�-[�������jZ�Xt��4�]��㣌,T|\Ye�*�ꋼ�1����C�G��@�î���Q� G��	��NUc��1���]fj91.��˨d)G�j�X�ڜ�[wP&���.��-�KE���A�q�)�ǄxD��	&�i��^�ݴ��ly�O�,�sK���!yka.is+TD1����a���2c��E��m��.m�ʋ�?H��^��-�n?N��J��h
�|�x6!��Kzs�?��z�D�����}�hlr�V����X 0�魷�ж=�X���v��$�{�K�w�KS��]y���������ْO��`��sqBX�:�d�
^��2ɚ`��A����hr|�S��o�B�7��Pa�n������&]3Y^wh�*��i��o�Ӆ
9Y�5 c�S��s/I	�(zS�<���)	[`�{,-Xc�r����b�e?J�>�z���tr�̎��.�,�^��
 Y d$ܳRo�,��p��.����ebIb8�V�ǟ|����G��x=�[�F"��J�� �` !ʯO��d��?9<Fﾷ�6��6��N�0�_ɥ5��0.$���
H�4�]e������I���~���;���O/�-ZNÓ:r�1�D�c2��pj��˦|1��݌ubl>f��^��r�w���;�0 �_��X�*2#.�$_���|�Yʲ)@����؉�6|�B�����KK#��of'
&�t:h�/ߡ��\A����+�}��H� &�n��iΡw�m�`�$�s)�F�'�`^��PRUq�g~�a@�2�x0��u��I��[輵�H�S���ڠ��	u,a�M��>޳u�A*7b����#qi����
Z�H��L��Z�������Y��E6'v�]���-�w�	9L�[K_t�Z��Ҽ�)�)���c���~:|l���Wq��	��P�EUb�|��2��p�C2�K��G�Jf�28<��˧w�b�e:�*Zɸ
�(Ϧ/�8�U����9��M/��v�RG�ϛ`�!��,_CY0R�qג��i`�_Z��g�}�:tl�1E�]�>�Ê���BI�I��\-�i�]zx��W������f�}���Q��#����-��ldB�+�]��CM�)��Mt>k�O~�n:�ܕ�r�� �/�������hbl��� �&�$��fԲA{�d!.��L��ū|Y�MM��ڦh������Uln���]J����lMPE����{� k��I��V I�.��^f��"웄�<Ӵ�Q6�����ڦ��4sƤ6���&��u|�F�V-c5C�l�!q�"�|�I�)v$e`���,�O�XMô�B�g�Z���ၔT�/�����y�h�,������)ӑ��)��ٚx���0`.�����Q�
���� ��E |6����+����������K¨�N�*-
iQ�?Z�W�
j]�
���V[�u��ED�P&��Ƞ�E�C�%/o����>�E1�k[x.�Zw%y������nJ�d3��n����s�!/��2�b�j�>���ԎAv�Ў\e� 4�g�#K����9ĺ#�(6ᾃ�I��P!iB15�Lĩ(51���3tZ��"����%S��L**w�o���^i���Ⱥ�[�;$j�tҡs/����$��#���w��j,�s��(@4��d�m���)x��T�cC�"4G����g1?����VHc<C4GŠ]�L>l2� �DoP��d�l��(ec(caPLRU�m1�>K6��Ҧ.��@c�	ˇ
���R?i���:���RҒ�HZu��AJa�ur�ĉ\�á纴��8`�ژ��<XP"T]M�:V؁�����X<"�E%إp��!E�w��0aJm�[C��ih�!�̑*P�kו�����+a7S&�(�R�W�s����!�,���ʋ�H��0��6�)�M��fٴ0c@ �A{ԷX�]a7�����2c�W�S��5A��]	�+&I��I0� /.��G��A�4��9�9��4����ąp:̡A[IF����Fʂ7�"����:���Ͻ�*c�`2^d<��G�l��gi�@ 6�o�m�
p�j�X����z���j�㺋��q��60K�]�1E��)*��	�X� �M�
��:����n� T+�".�yՈ� HǬ�̄�{����X�!f�Y.��
�,����@!\�N�H*������AN�D>�\@�����#�����P�hZ�2��D��Ds�� �,d��������[���8܉3ݢlM����
O#Q`���Mǁ!����IA�o$m�LZar^b���V�n��:Ds��?�
��)�f!q�Ͱ��ƟX���B��˧��0Q�by�Ȳr� $�̺�}��$lƪv�E�"k �M�a�f1)�2��#o�~�5�[��(ʾ�p;��x��R���2��L�d,2�� +�P�x�:�u8���Ĕ�V`�t��*��v�P�M�!��g�ƹ��AY�5׹�IK����3�3����I���y@�b����$n��<0�!;L�_�C��0/Yf�XI=�)��c1����P"��::*;�sı��c�%(��-fx�, kcy�/��	�e� �qrgX�E~�@��1	��t�k�u��ũ,g���6]	�҈%���Sq����-E�9���@���(�Ťa~�J\۪P����͌w	w��)C[⢔M�U�AL�b��0媋���$��gX[蜧��c�UT�:�� wm��J�eYa�d2+��� ����Ǳ�8VNQX��7�A�������b�����Q:l����F�e��j =_�U=c����Z*�Xl�a�Y�eP�6AĨ��,�,��CǄ:'�֓���@��v��z���suL	�s?Q��)�%��S�"'u���T��c���Fl�\�9ȱ2�Pp�&�+"�YO1������B�M�9n�2/"a�9a�9J[WZ�,o�zca��n���j���TR$�k4��i�q�t�ܳ9ʹ�|�@+�!6�J�]T'+A�h���הk-Hp���Ӊ�.'�졁��5�wK�2�G���ZB���8Tel/�[֌�ܴ�ց��̆O���D��0�4a]��p:�A�x�-$Rf6����#* 6JVf�S[A�!T;�0+q�X��صƼ]�a�k�4À�D�&��&BV`�����e٢+Q١���C`ɻ��0;��B�se�؟sDŻC>�����.��5J�zt1�8(�U�L݋N�Yp��M��\��d�8,8f5%�v7��L��X>�x ���(R*c���>��A�qEPZ���E���0\���<��ʳ&(vn��5�h���0>^`c�$��g�(PDQ6�'.N��V���\�pgD�3Mf���C<x��H����
,j�&h A�]�I�U�NVtLǶx�B(��D:��gT̝���\�)�4o$epb�����2�4{~2x!vV�І��@�"<PaL̰j yd�I`C�/�5�R��á��)VK��
��ayR�L�����Щ��@(�N,�����$�2�\P����T���A�v|xy �e&:���u�B%b�24�}��������7ޕ�c$�c
��[��x^�\..�GR��s�~��cQpf���d��p��'�ݘ2̨A�\�|��t{x�m[prnI"K��6���A�r�5���y�4�e"#��#l9�;�-���)�J�x��]�i2V��P@��R�}�6�L�Z����/K���-�i��)jC&����Π���m��Qjpnu�?��#x�4�Nw�P�Ia�DiP5-`��R�LG	�T��q��Z�`ٖI��'#�2�f�\б�����O�Bp�
,�M�$�	�piIj�?��h��e8X0��$����Bz*�-$�XU}g�Z�[�<vq�p�M�^��
�<�+�n��#|��Ǥɦ��`�	��`�l�M����:� G�$�%&�m
'���d��&=��a)uZTi2dH�R�{�����	������dHsJ�*i_}��m����%�ׇx��4�u)(H����$�I+WVD�S5g���ܾk�ƨ ����|C�s��������o�)J�H�L<�=��aYw�
���W��@0<td�x�Y/��M"�sZ�pa�7V-�7o>l��UW]1	^>nƂ��o�<&֔��c�vkF�q�l/�3lX�����R�ɲ���1�r��d���?<m��IpM��ۯ�QR�$�(�̰�D��l2��H5�/�����[�/������<1#�8��f�����q��Ç��^��Mh�l">P+���IQ�3��/��ڋ� ��z1gk!/�p����l��O����*g�O�����?�[�����F6[��+�&�$�/"yFy�XAY���E���$2�@Աº�⤋T&Y\]]�`��f���Jy}�[��P�
|�^�:�5��[���%qG����,��\H'�N���'���c-�4��x�7EEEؽ6
*:d�Z���a���t�kY^��Jy�X>E�8A�ܠ��ay�x�L�5-ñ�"7��IJ�b1�o8��<IO��q��1,/d-�4�<��g,0�4�����(U����2,�œ)� ��C<H,��l>�:3�aq3�L�du����v N4�=c�Ab�0����4M�$�0���\w҂E�Ѩ'����)������Ҥ���������qt�g���e!t�)+>�ݼiڞ����bY����i��yb,�,�Up���y3��9	&z�ЂF�򞱊���t��q�i{���`�w�G8���$mb|�#K�Ɏ�x����ph�qZ��䌜h�{��ի����np��izR�ǅYGl�ֻ,˞���T0װ3����ӹ8��q4�e�-
&��n<�����p�[n��FTxQ�,-O@\a� 0�u�cG�PK,ǛWh�����϶h{R�'�򞱐TUJ'9I��B��-�u��l��%l��C�u(Om�ޜC-�v����z��ׂ����@�����O�Xʈy7l���%���xZ�.(�MP��!�r8�F$�$��k�X��İ�R7�'��[6 e༬eq^m,fx��^BX�'hJ$o�$���@UҶ�?n8!�K�F6vI1���%l��놋}8ED�zb,�r�hSΰAzz�4�`�\��,Ii'�X'��@0�`�C˦tO�DC�����(��|4�Qja�ԫ@�P��2���tCJ�,�g��`,5N
��M�X��V�6�c��)���W�
�_��KaQ�e�tVa�;_�C=Q��`,9�ƆH����!qR@�΀6@%�Ib%	��(����0-dg�`�p^�'|ى��c	�da�5�'�7�e�65�2�!��������c�{szYÒ,Kpiahf�%�����IN�%3Ð�1A<���Ct�NjhBʛ*D�a"�Whgy�?eMQӈ����g�zpL򎹾�ED�۰$�7dۓ�l�fPWm��lb�P,x2��	| i0���͖"(*IYI�㪬7uk�g�q*��ߦ��
����.�h�
$������_��_v,��T�S�1���9��>U���]�.��VϹ�:;v�����!d�YUU�ڽ{��(���Eʃ�v�b5E;���N���K~������k�Z��"2�ݵwj���Z��$��Ҡh���ۗ>���9�Oc�Ѧj�S��p��͓�kMW�����a#�n����Z���;|�t�E��ܾ}{�����ɓ'�Ouuu����`�.]�駟��A��.++������_����«K������}s�M�o
��5��z.[yϯ^z����Qš'#�-c=��O�9�gU��ǚ갑*<�����^Ŧ�`նX���J�0i��wk�'��m��C��a��z�Y���6�6�2����ܗ����5���{�uۏ��3�<s�m��v��M�.�JI�z
�߿˸"�7o�}�֭gO�:��	&�o��}��l���߾Ohl"�E�t��Ui]qb�������7����o.��C�$��e�=�C�7��)�ٯ+��:MY'[��8S"dG}�!��ʶ��=��g%�k�W�[p�^�5��D"�D��-$b�R���*��7�ն<��r��޽?G5��COY�v��BnVM<�E��p�~
�P׬Y3޷����q�"nX;)�n�}Q�"T��;��)Hz6����D���7�^�:^˝�$��d�[����C�I��'�1i���>we�����C�~<v�����/��C-�[����^��cG���f��]���,�?	J�<�{S]v��n��5%��mߞ_-^�j�T$��^�~��7�k;r��gM~}��A�q0�u�]������uȐ!�˗//Y�p��/�����u뮺��[�J��Ǻ�U7�pUՊ�&��N���:r�s���5*F��)�\T6r���ff�ܡ�[',�����K闶#�۔��u ^{Q�OBXl�����D���Ƚwc	3pKo��X��n{0N�/�x>J��^��+/�V�ʕ�f֑����ξ��#��G���ohn*XS����� �����,\4�Q1� ���a�q�Y;v�og͚�0l�#F ��1c��,x\�4��𽧁�>g�k����A*����)������{��b�ͬ?Ʒk��Ҩ HM}<^;�X�.zf�������Nd�4^ح�+��ܰ�/x|�έa?��R=�&?�"kt��vw���<> �BM �K��<���9�X���͗�d����]5�X�����9Z�{O	�*.{�7>5{��򁱞�;w.2��w���2�L{�}ߑ�y{�̢��zpX8a36�1��R2c����������b$Q[7|�˥O������$��c����c�49������k9��FsCR�f\Ӥs4��⚌�ɵ�����":⡟]|�Xk�R�����o7b�Fٴ}��������54ԗ`ggӲx�B�c��cP()����P,����0�J�AJ�-��ƍ;�ZH�*���iih�k'l9I)���i����\*����-�3_������{���Z^���S�&ask�(���jb_H����4��$3vp~��^�#�v��?o���/�N7�ِ�$��Fk�Eẃuil�*��s}. �hѢ�ZH*cKaa���?#�|�ZJ�m����:s�����G�ϗ��� ��:5+��I8�;ƚ8ৱ�o[ǧ�=�~����?��=�s�wT�3mJ��LBDy�6Wr0j߮������)N�$#��?�?��|��kl{�$ca0^chw�N�b��eY�^={V�;|N(��y4�}�K�.��z=ƾ}�Vw���s�������s��Ds�����s�ҟ��O���K~�
ğ �C*.��{ܸZr�R�1R�H��k���%k*7L�������;�e*�����U�+V��éTH�j�y֑��{H�WY�X��x�IU�M��4_�.g�-uٶ�����ﭞ��b���c?[̧,��S��{�h��޿d�m��R)y޼yL�8�f�СG�U�r���\cg̘�^ "Rӽz�Z�E��"}z̏�}m�`-���y��iB����-��a�>=t`�[W����Ԡ��KW���s�[䤥�d�����.�]���Qip�Տ�.n{��b��UZ�ǎ̎C:���T�bѨ�Vr�g�ޫ��tK�9tC3M���VN|����H�r�/����k8J:H[.<��/�u�.<��ʝV�|c�a��i�J�xZE{ذa��f+��eYt���sJKK���k:uƒ9�}I�gn�,�ɆY���s�>;�_�Ѥ���t"��x�A���m��g��f��DS^2֨s.�=R6��􀑭��7k�I4K꒩"��Y�L�`_q陑.����Ā�S�<���JX5<�).fB�HI����Y����pF�ӻ�������q����3��,S_�z���i@屢�ֱŒ$%�ҏ~���V�j;��i��'�����W����|+��B��$���ϻ?:����7��Ly�XHS�����]�1�b݊fѺ �8��Fz`�^�v������_�lk�;���=Xcb�;�V��CZd�G�m��F[:�"�]}E[~�wPِ�C��p˸q;�ǭw�yg����/����0�G"��g�uֻ}��Y��Ͼ�aÆyMC&܋6��V�|s�S}��{����Z.�C��h�3�w:�׼KK�~�,^JNv�[�Bq3���Њ�[c^���Z���u�|��%�cI������(//'�K����������g��"�M�7�׌u�N^:�X��?B���G�c����?�2h�4o    IEND�B`�PK   w�X�w3.  )  /   images/b3ba8064-1e10-4daf-8b84-7882f41f3c09.png)��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[pU�y���s�IWo	��� �S�؞���#��y�8�L3N�4ɸM�N��#�8��8i�gܦq�&�qcL1�����0`H ����+�{u_�����+!�d�+<�t���Ϟ��������=V��6)̲X»$�T�+d �Kp�7ճ��t1����#��
9j�g�R�Ij�ӏz�G�Wh�+D�~�F��
�
�T�sAz/��v�f�����o�:�ƅ��\�h���aj�[�>���OSE�i\�A�6��utr��03^b�Ŧ��QLbm��n���kp0��5e�蘁�7����uuĸ�ֹ�!����9XR�1j�P��[͠��ZZ�itIp��=>�I�X!����T����=��`B�����&>Q���!S�ϚR��n�VK��1��=9`j%�����WV(C\$T�_�iD�}� S�9Ȯ�Jm� J9�1s���e�Ң�@ذ5��\�ˤ� A� M@P=l�Z�M�B�d^B�$��%H�4m@x1�P
&��/�F�N�	C��+�H�Y���f��I��BQ?D�x���$ݧ���iǙF�
y��蚗ka�J.��%�Gw��8�ؖGL^��n��χ۶[���O<�ܪ� x���(A�{��T`�=$U�x��T��a4Q= #0L�Y�x�f�A�1,UGZY����a6��a���ӶhƉhL2	>�H�$�X,���QMk O�4��Yԧ�c�TO�3�D��!mx3|�i;aZ5D#�,��f8J5P�Kwbn�+qO{	P`OG�5�w����k/�M�X�n>�կ����Qly����|����ӂ��Ѱ�&mӮ��Y-�ȨE�K1`����#o$R�t�$T���5s�Շ0� ��%HZ���qN^G�u菜C)ڋ#�Z ���V�Q�1f� ��Z��J�	6��\��Y��?��r�ӀaR���g9:�@�2��_�Ŵ�l����A�$̎� ����@8p��C��I�mǍ��:�̡�H,k��"��HH�M5؟��|(�V�R�vǞ��m{��W��L��q�8d7���q~|\xZ��D'T����V��ڠ�(N���$s�8Vnc�$���럔c<%^�u���)����h�,����������-�Oi�Xяg��NK�s��k��M�b��Z�&l���q�{]�M�����~$h���+U��x-D�\��m;\��L��mUM��Y�\�qhh�Q<���ю�Bቲ��eq���H��	M�$���<�F44�I4.]��$���������eGkN�Av}��7��Ň�~��@��c+�QmXlE)T ��!�΢7NGz
����cvhL�3Ez���m�v��፷��~n��c�*u�^�� gއ
�4ç.B�bv�E�._�N\Fu��
��\4� H(�������0��^w��$,\z�M
5�B��j��a)���#�{������g�{&Z�_!3=.[f��)�;���M�����P���6o��'"��ԗ$F�hy��:���]���/�z���sd�#�c0'�
��L,&�� !���@�k^Y�7��֊ h.��x>9�����<�XCćт����i�g4��uQ\`Ǟ�"���v���nBUm-�B�M9wQͳ�_n�P(��X��Ξ;�~��m�.�8?%��$�:���W�S}eT$3k�3�S?�x�ۮT Z�h59���  qCt!�HQ����7$���/n�!��qn8���ӄ3�c����=} a�x�����*R�U�$��d>^�O�:f�bCr���l�����XՋڼU��'6�4{��u	�7)���2z��oW	���%BX>z}��z�7�ϭ���w��-d�y<GY&P?�#gn�&��x�@͎3�"�Q��ߧM�Tf�&3�2g��^s�j�t��m����Z���H&�\��&�H`dd�`PӤ��Y�q� �W�1���pGk�5d\��A����a��l>ч�Q�g�6-��iž^Ы��L���[������s��e+5�a�(k���D��!�|S���?儑&�&*���H8�����۷k֬ѫ��p�Bl߾���X�lR���89K;�؅"�va��H1�|�
n�հ��=�w��k�{��vꇺR��A(�6?��[�jn��d�z �k�/��Í-ᙍ���x�ҫ	��}��;ެ�͋g�-Z�WIkk+������bΜ9X�r%�,Y��u�]wQn����p#��vqi�K��lF)\�	I^!y�S7��mX���o`�|A�<���x��A����a���x<a&3��;؉ža�M.�BY���؊N-=|9{�"�?x��W�k�.�z�ڄmذA��ѣ�����U�p��y}����p�tAaqv)��\�$?���5͓�'Ad�����Z��Y��I�7}���Vy�V�$�U*�l�S��M���Fg���x�5�(����Z4�ch5��SUX�h�e��%�k����?66��Q*��s�N�b���144�MW?.\����a�CFGG�T\}��>�eq���h|�N�ܴ���xЇ�m��&�X8=��um	��zEƚu��|E�]�H�u)�|�b��#M?�$��Ժi	r����x6�M�\g�%x��k�2�s�� 3���~`` �PH���i�����Ŧ��,ߍ[��a�#���΢����:ȇX�7X |1��K��B�L�IfU�^]V�J����ɵV��N�M��gSk�w��^9�a'=�|�X�B3��ٳhjj���l�[�Z����_!cca�B�*iRCR�O�7K����)dI86)C��Q�!�Oa�f>jcuؽ�9~�k���01h�u�����{k3a�����F�u�J��ˍ�`��ԷZ�=FB��x�}����.�����j�N�=�tq;I����t7������f�\oI��E� ʉO��ʕ�+y��(!�{�x�������PV�
������|�x���١,f�S���I��^�L����������[k�� ��dƏ��÷�dqa�5,���qV����g�� \��X���a���D'Դ����\wqo�>��l�I{:��%�埅P���.�:Y,[��<���7%M� j�����MD�*P=]�x%�A�VG(3�Uw܁�:�R��n�k���b����a��=�IN��1
����iFZo,��¨ac��ÞR�F��R��,N�i!��(�q?��	�9=�;�6�7�GC4�"	d��4F����M����f���.�c����J���:a����wMKX�5s��?��yUrY�b�8d�z!˩�$�!�\^';�9�u;�-j���f(<RV|N�L�^�]�	�5���#���� �w�R�'�*@Y���5���p��0�������e��&��Y.�͑�(E�:��������GQ��{:��$�h�ƹ�D�!Q�۲��Ѫ*�c8u� o�����_�ʞa`x1��f���:���\���\Vdƹ,���d�F f
/��h������E���mP�C�Y�8P�ͯr�zC���i����Z!���40�����>���R�oA��;Q�2SO����7:h�m.���x�p-�Ӡ,��`g�ˢ�:]zno��(�ˀ��	�Ȓ�sA>����q�NS5u�w��ށ�ɠÓ�$a�Nb�*Tuqs�����&7\5=R��\����0�̗u�
Q�`�uܩ�q.Kȷ��Lg�ު8:�8�C�pL[����M��	�/b�ʃ�Խe
{Kt�t�6�Ǳ��]��ea��8�m�r�^E��<�hvB ��8q����Ny��!o�PH� ����iE�_�J`�/��߃�'	d�l�ǻ�B:���]}�!�Y�9�9r���b����C:��&�Py�f[��f��rq�4~C�����5���1�\�;�0�:%z��t5�
������1�:�l1�&D���@��ýi�������L<�@0�]*yy,��G�WC�(������X-��9E���^a�t���]j�m�9����,i���;k[MHg~�OB5,��7७[��
�B2�o�@��S�P�L�2i�0������p�|HAy۹�_
g{��Ÿ���/ۻ-eb[_V��磣��P�}�e2#U�����,��?����� �k�y���oߟ���Õ�,6Y�)0����x+�g�?"��,�qqy���Cs�
ޑg���@�NazNS�\�H��KF��-Ӳ&�ej�������x-�L{�0�[>�b�ie���
S�'�?�Pz/D���Z*nmdu�̠7�:Za���#XAÒ���yf��K���,Р���=�gz�$��S	��*
QГ,P|��*�'�FN���9��ȢF��{9����FOnH��W>ԫ*����h���
��F�j���ZzG�z���Em��4�!��4�]sE�5D%�1z'��q�F��8ˑ#�Л��T�4�O�X����\[��b�u�ҥ��ə������Q\�
��W�~��'y��eW靲J>�K�X�;Ļp����a�gހ6Ta��=��>|޼	b�� ���G�e�%�|�݇?1Vb�h�u/�|�hy�ߓ{QO��1އ���Qw�˱B��W�4N�A|ڸ#��1w/�>�-ح:�|�R?����Q͟��UE|��-�K�Z��AuO������[�eA+.�d�D�(I�`s<���e�ڟ���*��������~�����l����~�};���1������+3�'
ٳ��Z�j�:��*�A�݁P3o�P�v�l;����10��G+�N�,� {��lP��iō\K�a��3e�7C�VzW��ho��#S)��䯁�Q��t��63�@���MR{+̆�1�d6�(�pM���d!b�g�������9̭���s�t"1��2���1d�΄vA����F��a�jꚚ���b�R?�E�*Y�-��7v��v��>,��W�)l/���%��P��I�е>+�	�b�!aI��߉���6���A����;��N�[DkS_��������+���'��lwQ����������}@��3~�[�.BYF�{��y�ǲ|>���F���vr���,b
/�w:o���2\犄�$����N��i#��Ϙ����ky�<�v��ौ���$�ARb�|-W�V�p�@?ѝ.d���D��	r�~*��DG�����j�����!��)C�X*����΂wV��\p\�9;�KT�LJ�X�sd��%	clݗ ^�.��я<^��t�p�هwm*���7����m _���!�D������,*?��?�=�m����O������y���e&3���x�b?;G	=�z�p۶�w��_$�~y�|_����Í_��aN��o�6ɩ��s�w�?wX� {��p��B8�����Bj�f��b    IEND�B`�PK   �u�X.D��N �M /   images/bb8b4d0b-321c-4695-852a-55709d7923fe.png @@���PNG

   IHDR   �     ;��   sRGB ���    IDATx^Խw�\W�-�n�\��9��j�rN�������`��8�`H3�G00�q 8��s�d[V���S�X9��{k�*���ޟ��>}����u�9����k�V���p]WS�����/�@yP��p��몫VAmjک����e�lջ��ܛO�#�)c b��&Q�����ôl7TȪ��OT��W�@�4tM1G
�,�)���EM�,��uM�#��KJ��)�^R̲������@ST�Q�R��c�m���-��j��+��p�K^?�Hs����{�)JY�hpm�*�KW�r��Wo0Ӏ�e7��>�P}�G3\G��N(l�����z����r����ݏ�z]����\,_���Ǵ
V�)�ڀ�h#�eem�l9e�q��*�b�E�lY*L׆�±Wu]KQ��9TWq۵ǱU�qt�,k����~�q�vt��*\^���P��]�>\> ^Gq��
�[���X ������ .��N� ��؊m:���xT�Qt��g��
_���J?���UE�{�8�⸎��[G3ߧ�P]W�!Ô���
��SWuશ���E�!:.x�2n�Ǡ�Y�w?�[ރ������*.f;pm۶����	�*w�.��#����Y��*28��F���+e���0u�p|���=�-�����^��3_��Uɿ����a-���/B�����r(�J�4t�e��A�ۧ�MN�bk�m[saۜ
6��3丰iG�b�PhT|�P�(ނɝɽ�b8��	��3^y�u.�a�
D�����E�"V|��h�����*�Ů,���{��4yO�}|��︼�7.�������?s��w��
E���~����N�����%�Q����2.�Q�i��h��m��T�J?&�ͻ�^�Wo�\%e�~~Z?��P|*\łj8PT����CWB��\����o}��׆5��o~
��;�.��7 ȕ�t�ꃪ�a96,ג��E��@U`:&���E��tE�|Oٶ��'�����1���H�(�\Յ��Py��*�$nC�+{�q�ٻ�gl�������voBu�Mc\��s��-�7�7�~V4M&�����-Ck���Ò��F��������ާN��͕���υ��gr�C�U��bht9ޭ�������7&~�c���x�P�/�*���*st�r	�h��/����CP]��P���;.���׼�O��O}k��f�:��̯�Wu.�z,�@��`+>�5d�]%���hP\��z7Q� ��F�}�	14��K��lۂiZ0m��ϻ� "���qm86�{����jr�ғ��\`N�<�3,Nn��8qܻ^0���"rs�t1۴��S4U�ŀh�P�IW
�J;n���AϪ����g��/�_ަ�,�L�G�^#�b�/�OxޥjX�����Q����-�獟�#��b�g�jȮ�T�ƬҎt��`:
LK���&l�N� ¿�hA_F1q��7|��\{B����C/�����,�*t����y�v.L@�`�>X0�8>q����딠�TG�ω����W<�q-Yx>��}:��M�V��Kc�?N�eY�B@5Vã,�Fo��İY��i�=�ޡ���cT<�x������d�+!�Cu�b24q'>$�V�j��/�x�=��BvVé,��P(&��r� ��`]9��7:W��*���ÂK��l�дx��p�~hzP<����:J�#Qǲ0�|���X�`+�{�i�n��'>����uq ����x���K�`����d"0��i��AB�N���*�,�0M�E���`B��r��{1ޒ��B�`:�	x����4M�|GTZ��	��z��zᰂ�*����'N�����L�9fU�P�$^�|����W	��=�:f��{S�
�*�E�����M�|��2���{c(�=,'��X���:bpm}���H�M���,�a�%X�#kcZ
J�[@1���D�D(��H!�~+�͙sn���W����Uʺ�j�����ϯ���4\=�-�
El�N|c���+��T��G)=�P@G0�O�ñ�J��V���0|(����kP5��)\	eUU=��jH��Í�tR`B8��<�D�ߋ�d���ǀ�౐s�d3T��D�.��,b+zX�x(��=9^z	I�d�&�@o�Dh��Q�mZ%xJlZ��4f�%�웋N��&|*����F��\��8 �2Ũ�V>'�/���|�F&o��$�X��U�\'�0�P ��!'�{��n��MW��<��㋷���wz��[���n"0`[z\��F̡�
�f���.C��uQ���LR$A(A ������(lYT_6�Z �?�"3&zo ����(��C��7��ty�d�Ъ�Z�9��%4 ���J,T<�Jl��D��ӽI��	r�KU��D�\�D|��@�(�,ج�-Z�*��tPe�fއ�g�C=��a�JV9a5�P�H�*#G	!��e�45?tAJe��hi�Ǣ�31��S��$���t�r���cמغm7�����H"���CF%R�"�i#5�������)����-�_�w�U}��<���~�k��bG����+irc�l�]�_�0�l�P˖.ĢE���5����(�
AO� ֭ߌu����A�Զ#�G:W��B�<�7����.��&�щ��8���S�*���x�ޛ`�JXa�_}����h`qԉ�K���C ��*�^�j��1�|�� ��V0�ê�u�Ұ&�?1�����U�"�>�k"���Y(N>�����1kZ'��N��"TC����ЁT��Ν�e�.���M􏥑55��A�SP��[�P�o@/����n���|����ӿ<~��O����,��b���B���@PC��DmT�E��Ι�\y.����f�2d2){���H�h-
E��������� k�K�PU�P|O���x#ӱ�q,��������D�êz�
h�~�a��&e�t|�ߋ�d�}WV��1��FTI��4�������z�f�����=:E�W��M�K�00.b~E*�@Smz���ҋ�C21�TDMM
墄eM5�֢���
<��+x��ױ�o��|�F��9+*��q�B:��H�N���[?��bXz��G�~��9Xn ��ç�*i6ɳ<�a��X@���g�ګ�����0>:���1�P$�`ȏB!'�16�FCS+:����p
���O��'�k�b��GIB�n愇B!1f���_������]�jh�h��z���\�	�U�gYCx�u��f\�
�Nê��{.ǏU��c�F���߉�[zAhnD���҉��bQ��|buQ7_�\q��0�Y�"
J�`��1���0C�Pt�xÇUomēϯ����QV"(! �0�E�J���N�}�7?u�'�X����>��k��/����4�.�/֑���)3?�SOZ���F4�ƑO!1:�GX�\8�	��/�Z6���L�-����x��klG���<��q�F_s�5���T��[�Y�U�+���S^	<���oQ�|�S:>1�a3�
X��M�#2�I�Ta����cۡ⵪ia5y�%��I����fO%�ⱪ �����*d1\�C*�R(����V��7^����@�`e^�P(��r��e�!ke;�$Z-�&a<W�s���CO��=�(�~�b��EBF�����-�r��>s��'4�_��ׯ���U�ٗ0Q,�pLW�sP�Ž��<����SZp�uĜ�.�F(˒%0�)�2x��ǲQ*�D��?GM]3֬ߌ�����}d��6����� �7, ��Ya�e~I	T�E�# =��f��DC���	\�1
�9�{=�q�:^��������d�Qeԏ3��-LJ,�k�(�J����<i`(�OXJFރ���:�v1��Xq?PH�a�.��������n��(��b�\$�*��3�����d�[��n������Ϯ�P�B��	�x~z,s���˧}�z���y�|�͟�P4u&i�*�r�`������W^���)�z��-0w�HiX
�����k4?�%�����w��_?����S��waR�l/��*��
�2'���H��٫ \B܄5�h�7��j2p� �c�ci��5o,�T�~ǿ@x�J��]��
��܏���Rx�*S_��`�=f5�Vy����{�ڨU�j���碜��o�W_v&�?�`��Y���lz�1`Sۂ՘]��2�Z'I���ڝ��]�c��~h��������H���B�/�����n��z�],�����g�5ʈ-��|�ʗ?��]���f�����|N�(���bQ�,oZW��y��U&wʌx쩧����{���1o��N��i��H��;,r�c%)�E>����E����P���
��e����R����S�Ŏ��JiJF�B�GJfك���EhHn=Ò{`��SJT,�x�1�Se�e�L�%������%���WZ��Z&����A�a��d��}͵�F,B6��/��!���z��4��&E���@>�F$�GѲ��э}G��;������4�6�"��)��_u����מ�n��o���Kol�����^�uh���߀�Ck]@�k�����׾���A!@9a4�#&���,k;�P\Ky�ca��"ʎ����رw/��?�m{�4{	��8�${����#�C��I��RÈ(`	��~�C$d�
�Y*�|Q!+�f�(��9.թp]U��{�`Y�}�G�����(yEh�d]Rՠ�=�^x9��΅��h�_iU�.�O<�4�\&�"���(���
ou�I���� b\�B	!�AD��JԘ=���߀┐�¹5��GJ�2|���`��}�i4�
A�8�$k�4������j���<��md� [�"��VN���)���|��K:Ս�_�����|�G�������~�3�� BJ��\u��H��"�L
!�KbX�`	�y�}�THpJl�%���)ƭ��V�ݏ�y'���ޣ6Xt�ީdq�������x��V����P,�^)�U+X�|R�ق�~�.�pb�&�r�SY���)J���~ =�W�4<���¯�M2M�HX��e��%&�x�|�$�� ��\���gh��r��^	��m�(���$�J7ȽqӘ6�>�����0�=m~���Pl�s &��U��eKe��Z.+ ^���������?��~<��ZgU�4v��A��+N���o|�W'8\V_��mw}����ޑ�\�hQ��a��D]HA[m 7\{�:�d�9(�>���1H��TA�C)	=�݋�|FQNzsKF���{?Ū7��s�r�����~�cګتJ$R9A�Mp�̑�Av��1�|ƅ�g�g�xM�6Q.�aKRS�bh4#ʂ��ҫ���
����{���ǖ�O��¯mc||���*B�y��0�G�Q����P���ɐ��|� 4#�����F���]�0�?��{ueR"�b��BwM���,2�{q�)�_��:���i�4�@H65eG�.,��S������Zq����MAm}������}O��d�@k�L�F~77r�������|���}�g�]��GG�S�%�}pK)��fLn�u�+�/A���EP��)�)�Ix�[.�&
�LO�P*��Q�LM-���ĭ��	��ރ�'�&G�,�R<o�ɐBc�Aq�!��*��(�!�vŅv��|�⠔K�\����bDqM�-���hoCc}����x��������ba����PЄK�-O��	,��n��i [,"�-B��Q�E�Q�30��$��9����8�ezo���0+�;zD1�
�*!q�b��<��@1 `r�dՇ]${wc��F���߃��A��d�����;hhmw�"��:�����CcK;��㻿�~�98�8�'uVS���KO�z��?�'4����ޫ�|��_εz��!�ⳳ�j���k���'�C9��U*�@�A���E�9�K�#
 <WK��8#_41u�t��u'��?Ů���]�hMLnޡA�h�؉���ra�6�Vv���A�M�2I��9������&����;'���	������ש����^镐B�����%#���}���齚��ߏ\6�T*�|��w�b�T�Lers�ꛛa�BH��H�3��Ǿ}ؾ�鼍"9;R7�
�p���vŻ��No��?���D�TDH)#pP;�ڠ�_��{��\+���r�(��J�-�l��K�ĸw4;6(�P�����~�xn�D����C$�a��.^>��o��gNhX���ѕ>���e;iX��H���RF>ُ�(.>�4|�򕰋�
Y�KC��;�+�T����,b3�(����D�9�>�����P�7�}�\�"a�R���%�z�`��C�z���Q�z�BF��OU1����M��fLnk¤��#Aف�V�P 5ш�l�]o��N��H�K�Ī��uTccc��:������1��jlh@m]��ca���C�cO&1<:���ಆ�F466�,%�W�u���s��G"���`�P5�}���1�䢋���4�%�2��
�� �#G�?��y|���n��$Kc��>�U�̫	�Fg`�,m�����ϭz��ѯph �Ǝ���~)��l��E7}����??y�_�x���ù���rWj&r�����ܩ��§nF�pP̥e��l�d�=骧��HC�PS(��>4���X����}�y�OY����P	���� �M��BX�E١A�.�V�,�,�`���"��h��y�j_	!4P�H(oii�k���p�������8z�(҉$��	������9�#k�A�Ecfq�y\F���$�a��niiAW�tvv"^_'��	�3�H�H�QU��F�q����[xs�.�����%�Eja�Vl�`�A��H5�/�4���з'N?i>���/��6�DrT<��.)����C����T(,d�K�,#����E׏�v7�}�Xz���!�DCp�c��L��_��'4�;�}�?=���GF
�X2O��%�v~7���|��k�h�t���k[D͢�8E��"8e|,�pMu��ذe+~�_?���14v/B��e*�6t# ����u��l;)�V��ʧ�+�>m
������������Pu�0��Q��	ط��}�bL��޲Be���BJ[�@�?@,��+�xXCFȫ�@�Ϟ��L8Hfs�
�9��t�XT�-���{*�_��sf���M��\߲���w��h"�Ǝ)h�:�/���`��mxcݻҰ��w�Y��z���j"c�)���ac|�0
�A|��u�
��8�GG
�
�&#E�{�����`��L�D,Z���<����W+2���(:�u5��G`���+�ϸ���O��z䜇�^u���´���R}(���<��"~�8	7\{B~��Q�e[
�$ߊ�.��ᄋGr�^�F��ځ��{���ށU��D����i2�������@%��X��9(v������9�8�E��݉��������ȥRxs��X���=�|6'��H�j
G$;%�V��J7+=D����傌K4�+);�A�N�*B"һ2�0�"����Oc���E�TFM]�Z���=�����ٳ0{�lO�fH��c���K��j�Z�1u�Re���M���&��P��-�(�.��(�{�J�-5��ֆ�|
��v���7�����\�bdx@ԥ+7BM,���]�\���@[{9}��z=~w�ز�6��crd t�� ��X���]7~�������s~��?�ul��6���f~P�U���׾�r	K��!$�F�T�̊;VB�dWT�����D�8�7��z�)M    IDATO=�9^L�>E5�l�㾂��gLVY��>�F65�X؇S����@פ�}
j�!��c��%�ض[6m����0��'�&�PNJ���V)�+�(�EC�s�br6��FF��h�h����ڷ�*�'F�� J�G�c3IR6MH�� �"���$i����2
�2�%S�z���z\p�yX�p>�Ϛ!s`f�8�s����x
-]�:g!r��_߀���OonC6o�uH�`��S���P�[����"�����W���+ܖ|7�? kF
�����de<��s���E�h	E5
%�
�I���!�x�;Փ�x٬���>ub�u�Cg?�ԫw�v3�Z�gXL�)S-�ƊȍbRs=.]yNZ2s�u�T�`l,�\��Kh�\(h��(�ݶ��!�ۼz �x]3l-G�TN&�@,@���.g�M�6�����'cƔ��Ut�� ��-[�z�j�_��R�q�#�`��f�2K(�q��S�{me䯤�Sj��0�LV�%�B��A���xS���ʰ�)y��E�<E�O�/����1#�KJ�`PBr2�A�hʂ._�g��sfτ�q�1<<���b`4���)�9o	�[v��O��]���D��Z����x���(g��ȍ�S��k��I� �>��H�J�`�ĥ����6<���x���� T���V�%Ő��0�T�%�7~��İn��ɳ|�;���O+)8jK ����%(Na�A&9�,�Yq�<,_�-�m�ʖ-�T�B����~��n��>:_$�`$E�� �/	����b#�A},�%�f`���X�`�0sj'� �z�5<���8���lz#��|����,��}K-M�,4�j�x����w
��<�ٌP��y�Oz �p� �b4��a���T2�\.�������35╆���O�?'��PP0-�M�b	V��p0��sf�ܳ��ҥKaĢ�{z��i�v�&Ә6{�Ϟ�t���|o�s{���B��4G�f>�SBzl ��Cįa�N�yƩ��Q�F����a��Cر}7�������Mp|5�+~��8��_+#���/��;_���Y�~��{z����� q�D�墸X�z��'FG`(��q��ڌ��.��O�I&�k�m>|�w����(J�b�t�X-E�="E�AX8w*ϛ�y3���T���m�]�e�z<��c8�?B�0Q�u��qL�������4uXV�!�`?�q4�`m�;ﴷ���l�F9I�/��wT�Լp*������nttC��$�e�q�(�H��b��x��}���jj0�Hc<�A>_��@�P,�fL��SO�i+V��c��hG��֭�%�]�x1:��������Ko`ûېΖ�+�0ˎtIX9a�q>	+��$��	c�\D,�,���6ؗ���A��ʖ�Z�]y*U�<���!PܠFR-������G=a(���ז�����z{����Ѱ��/�>�K�^a�f�H'F��9(�)x� ��pB`��Y+���jz�f�>�Pl��0�tMnǩ��ӖaRS-�~p?�{s5�X��ݏ�HT<��mI�W|v��1%���˶t��A�DwO�����'O�ܹs1g�\455�����N�ou��f4&���jÄ�U=�D�#X��^o^��)�<�E6�e��Ç��{��8�\�BV�����92:�d&�u3:r�4�,^��\r��uK���tdd��Y�P�KN;�x����S/�®��Hd��ґ����P���.�-�G�$�Ơ���&�/"�A,������Ï���L��B�v`Y���.����.X�}�w����OhX�>�������o�8��T�p���^)�b#���S�cq�V�����k�^��M�	�$�p�s��bq١��`@C,P��p�%+1��N���_����x�'p��>4���'����̬��G��ދ,=��D&#�r��N}��gbj�4�[0_~���1��+u�b!_�v^����I�����G0S%L�А�KC�����
&��=^�l	���\s9���b߾}
��L	����H��/� );��Y�T��9�p�ޏ�3<�9�7֬��1u*&O[��T	y�y��z
�������$ۖV1�=F�Jy�:RXP��1J��c���2�(��TTX�r�8�V*}�)�o��?��?�X����cw����"G��т���R�'�e��{�����}���L*��E~�A��p($��X �(B��BLJy�M��^}��8��˅<ʙ�nڌ�o�E<��-�q�P�F��>OJ��R&��qCa�uv`�i+�줓oh���#�ϡP6���#G㢄�!�.p�����b��.�|b��R���碁�s����~?,fX���� �-�"����4߱3HlܹG����1�&�)�<�����iT��oļq��+��܌P؏;�Ɔ���6O:NЏ����_~
�C	i�Q}>�39)��P9�l� !V�2��F�pe8��_�Y�fњR�$�%��Q/�eV�2�����zb��؋��y������[D�e+j1)Kc�k�Z��j+�t���z�.��X<f}P%d�5��c���5,]:�\t��.� W?�ك�|Zxڔ.u�A~+/�1�ҹb�h�hLąL��� �M����?_HH-Fzt��Ò�W�8. �`U:\[[#��j?��=5�Va�ӞT�gMT6N����76��L��j8�7%=�����E���b��s�Q`b��H������+���>44 �&J���
��\�ꐋ.�_z1Ԁ��!�ر}��X�l�gvb�$���3X�qJ��<;�?�E��q�)
��"�5��Q�
�"���rv�1� 	!�L�g/:��S?��-��S���#�ܹmw�������c��ɵ�������rOo��X[I�E�P�j���)���X�RӦ4a񂙸��s�O�"=6�Lb{v����0Z����^|����K��
崛��QY���V�u��8��h�4	f���G��Ho��|z
��4(d!M�>�B__�`���8p@�����蛙�z���L6-���4Nx4��o�y��`����>�[�_MM�x�j�H�4X�e�D�X�r�X���E��hZ��e\���Ƒ#�P���`hD���)x��5`�Ÿ���Q�P�T2��w��o �͓�`�)�4௏����=��TIdŅ=`P >�7��i��.E���9ej�t]朸Y�>T<�g##�L�e/X:��?����=�a�����~��;v�8�K*bH�j���׺Ms~G����D�A��)B��@wY�rq��sq��Kp����4��9�l��&�U��4��0DC!�c��H<Z;&��s����K������ ��چz��5^�&���ڵkqp�Y8�z���3<P�P߄p�e�	��\F��H�䤳��vtt］���&�!�،s@o8c�̟?_�輹s+�!�z4j�T5���3y��I�BO���O`hx c�	���4���^�8����م}�z�[8_��{����͛��`��%��5��u�H�]�P�Z���2UhR�e�4����0D^�
���oH�ұ��W�h�H�T���'_�ğOhX~��y�������?�oK
����h�l����D;e��3i���Gf|P'?���PFߑCȥ���s�c"P9�Ch�R�X�+	K��
hlj�y+/���]*�o����GG�3M�-���0�c8t�V�Z�6�����p��.��g����*��u�\�$�^.S?���;Y�v�3�j�,.^S'!%96.�κ"���Ja����k��JBap\]]]�5k�d��cⵘ�UN	d���ey_c[���R&#�߶m��~�fc�q���
f2Ԁx�K��篼Z@G�`/֭_WW�O���ï~{I!mG*�J6T�Y.հ<��;��h���kIq��DԨyYdհ�����:>��_���'�XO�:����;{�(�A	���a_y�����*�����Į^=�Y�D?fO��_�>�Dسu+�:�H �|2�0�������S*��#bd|�P@ ��W^��I8|�0>$�P˅o P�ū���Kxꩧ�}�N�C~�~����+q�I'Ix��!.�岰��!h��XW�w�Qѫ44�y*��LYv��,0 �g*��tm{�@z���u���o͚5ؽ{�������'�,*�Ky��<Fo������B��y��޽{��ؽs7���(�Eq�'?�9��A���o\�C�c�%X��4���0����8p8%��i��f���VIN@��4V|>Xf�cUd5��`�=��d��:?�/}��'4��}y���=�����=���Q1,����~��N)���ܖM�y��[F9;��������-AH���O!3>�cAD����fYR�#Hw5ea�Kh�.��.A&����;���YLN<�A��C�����Z%��sΑ��`�"YH�%�ᄋ���Ѱ_~|<)a��Df\k��P����Zb����4B���dѝ��k�M�@td���?ϰƐ��~$c�)�=�\9��^����Li��m���"$gs���/�4�A� ���������}�^�H$�t&��7`pp��]8�q���_���x{�Q�]?�G7P�J��Zl\����o�d�J���0VM8�H8�r�������+��?5���y�����;����y,�	�E�X�\�E<�'��\XVٙ!�<,$?��fcJk->r�e���xk�K(d��BR�SY�������@�
�4⍍8��Xq��D�8t�06n~[�xS:��y�B��f5{�1�WK�-Ź�'$hcK�`+�h<]�h��^�����Oג0�	����FU�"�ez@5A�\��Z ;�=0OH�Vտ�fU@�p�5y𻪽���K�W�¶��J�@]��,Y�X<^!�fᒈݚPW_/�:�S����b�w@�h���Y眉�߷-�R;$�w�!�N�Ɗ����#)��Ď�H�A���T��Q�ʶ�wO�S���3�j�X(�p(�r�Ͼxy����>���/Ϲ��'o{{W�y���y���ҰH9T���aI{���ǲ�R�#������/�"��>��Ckst��8uO.��[Md7d����KK����*e���}���j�{�4���ׯ���ߏ#�	P��5������O�Ԡ^&�E���������%؜I6�{r���xD�d�YL횂t6%\��,'�
y���H8�\X������r��$i���q$��f�BW0�Ҡ��[�7nƮ�{0�{�:�l45���Lf���(����"��ql��c�ƍ�Je�ܽ���*(j/��b4��
��a��?tS���¥Kq���y�y��q7�.�+\9K���k@�xK`�jK�E�1
��Q�u/\��՟��ɟ�а~�Y�>���_߸g��G���E8�_Կ�
9�a|~]p��`("hMȇ|jN)�����K/@>9��xM��&(&uL���D,��~�%���514��K�Grs��w�n�&Y��
��a�z�{�ط� .��b���Wc��i2�@#c�ӣ�1 .��5M��Y��Q.B�S���>4��c��
V��#��9IԔ�"�l�*���Eb4!)Ho]9�N�fIj�^g����^J���ՌP�*�hJ�Y�ڸn��X��%D2�d�"�뎧hkoA[[;̊���5���~�� ݐO"�)���I���;m߽�6mY3�b�
�'���=���U���a9&�#��5G���$S�1
0x���HAM(���!�������g����Wg>�ȋ?]�q�����F%�0�sHmS$)�dة��Osa����c��)����3x��Q#���"H,�V�k��aԠ��~,;�T)��a,���w�"A��/�];w���\}��v"_*���=�����_�I�-�P�G�;�����Wh������G:�����C �k��1�W�D
��=�X8$����H7��=�kʔ)"?�7�6���+h�4.�Ħ�	��$۴�heaŏ���zbٲe⑉e��ƒ�2~6�̙3GX|��߽���B	C�O�102�����O|\�b����oaϮmX0�-;{�˸��'�«k�h5P}up�����(I��cD7Oâ׎j�:��'�����NhX�>���{{��ol�{�W�����M�Ov��2�VNlg�e#�3�(�I`��N\��K�\��u� "��d��LN��f\lL�����uL�"*�d6���Q����c�d�n��v�>���b��R�܅�����Z'.P(��#�	�Zhhcc#"�,\4��앾��I��־�^`ɒe��k׾!�������`/�7z�����Q�u1,�3���Z��@�0����G���1��T5Tx�$K^Oc8*�(�K�i��x����{� ���j	��#C��H�P�2}�l|~2i9**�t*�����A����p:�LA}S�W�~���A��y�u�Yxw� �{�Yl|{/2%%ǀ���T��o���(�"��H��E�'}�o�{'6��_�q����M{�,�/�z,!;���!��12������.@1=���q�uW�ʎ��'�����
�l�e���Y�s�?\r$��<O"sn���a��i⁞y�Y���K�:u*>�яb�ȥ�	�#�6+�
K$1}�t��w@���v�V�£�>��o�Y����3�bQ,�;O8���1��O;]0�`� f͙-�;�E>�EK[3jk����C(yqb,���Ai�hnn����o7��Cԡ�g��c9����|B��h�t�+�T:fh��P����9�D���;o�,_&~z=�A�`(&!
������X��-�,��z���/�r����_/��r�uo�!�7s�)X�t1^]�w��f1��Q�O2Q��/}�%p�ʍ0=V0���~\���[�}��'6��^\7�O>~��-�W��/$M�rԳS�}�+]��t
55qhv	��^i=���>�-�G�*:�����X(,��J�K�+�t�gCCC��s>ؽ�İ�䓑H&�K�ܵ�f��g?�Y��FF��OL�Ѐ�1�����n�֭����*�s�n��3gΔש8hni��f �C*��F/3"Jr2���/y"�}����(�:ڤ�י���u"ʣGd��?�z�@�͛'��;�#t��%X��$�	���"�180,?s��rU�3���
��Q9�hАv�ޅI����+���%).3,O`�E�^z	���yO&�w�A�L+W�ĥ�\&<�-`Ӗ�ؼu.���hh������<���,�Y�/�	xg����%x��K۾��o}�'�Xϼ�~Ɲ�?��uo� �CA�a9���%<�]�d��5��1Ĵ,>����&ּ�J�q4Մ���)r��9W<q��6�Ț:��x}���锰�S�����6o�/� ���O?�\r��7b%���&lv}��h8+W�O�m�wkk�t�݋��{�*��SO>IvߪW_/Hp�H��Ȝ�=S&wJ����N�lG[K3�z���Z�f�M'SR����*��14r�ɐO�:E2�ށA���P����ċ�VY�'���"��V����]�њ���4�H��[>)�mxlTB%=3=WM��b��|[6oDmmT67��� >r�G�x�"qܷ[�y��c����#�Ҁ;�{���C��Xz�/&ԓ�6?��I�4�CM,���!�3����/~�����kkg����~���C�MUt���Q�bA�}��lVn:�ɢ�������g����y��z3�&�%�S�� �rA�m���/ �XM|����R��J\���ױn��u�9������$�L���k||S�uc۶�R�8���er��G�d������kV��?w�x�Tr�W�Cڲe�����F�V9tX��J-o1�\!'!�m\�i8x� A@��mm�G��    IDAT"��S�JH������-����ӲI��ldxL*�lU� �7q,�E����{��!����x;��믿�j�!��l�𡵕�����lz;����38��t��`΂%pM=�I٫a�$�~�E�3f����zz5�-3`�[�a���	%m�ш��?��qμ���_��	��՛g�q�ÿݰ��Yi4$�����&�|:�xM*O.�!ݼi���g?��k^³O>���Lii��
��O�,�4z?�ı?�tu4�t�t�`���%���ػw.��2�{�����,�A��Ԟ=���6i�$������ŋq�Yg�'��]?g���54(rWlL%�Z��b�&��� ���q����F�%�m���X]�����b��`�CK����#�#OE�ZU7�癳���ٳWd���f`��S�m�v��� 0Q�=RE���k0T�p��64
�B0�!��6����w���`%����FM���M��;n�`�Q46�K��h���?t���5orc���u������o<����s�E;a�q�h+�TJ���gOt�G��9���������Ϯ�󗇞���v�aRV��T:fI
&��+�TR#0�<���_An�0���m�	�1c�T�����u�S_(gU}�0�<���E���u#�$f̙!���^���.�y�'���^��4M�04����+���mܴ	���5�;�m���1�[�3�֦f,X8O01
�sb3.>K*���!���/Ac�g�"�`�dur�\�m���ر�{˦hii����I�m�I�<c�l>e<�����0m�L�ٻ�<���I���X�Ḉ���x���:ሧ�%>�����}�qL�~��O"����˦tM����?��;��KᝆJ�\�`��ȇkl�o���^}�%|�ӟFیY��o���Q���Ht9S�2������J�bYw��������֓�o�{�}O���-{VXi>Z��ݢ�:�j>�Bvl v)�/�&t���Ϸ߆|rs�MG]$�Ȟ@:���&A�܂�d��φQ�w��hnm�c�xk�:q��\s�����p8�\hb$���
�NP{�i���܋��f\x�y�N ��i�,��~��5�EN���9�\��˗�B���HV��b25.N�/
R�@o��@�بX��Hw�-���(r��)
T���O�8��<f��1<|�G�g�y*ּ�vn�*uɖ�6�Hof���� �0:<(��^K�U�3���=^Q���n�,�㤁rNn�çc˦�x��'�ͤ�t�"�	���)g���/��Dr �U/��ޞ�����#>���������QP�P3��V	-�qDI���i��~r�O��o'�X/��s����w���u��A�������;���Ǌes��ƋO?�7_}3�:���$�[2�Պ���~�eR�c���QJ�'wtJid�ַ�?��+��N�e
.6a8� �K�'	�������6lX���8�#�"�e��[k�b||3���.?|���뮻N�,�4"z��_;w�D�6&��顣��_�X�v�B&�Ŕ)]�1�D���"���kr��4���4\���'��O�O��k�41����ªW�ż��q�+1::.z+~�FJ:�ܘ���#�A�tNő#=bd�-��� ~�Qy����%�ir�E|� �twU�v����ȦS%h����ӟĴ�s�����.֭}��;q�Eb�����߇�G�pH缺p}MDHqd�tj��w��_>�a��ڦY����;ֽ�o����fBv6���s9��D4���g1ڷ��ט�T���6)B�� �4�퍥R�<a���R6���t��{�ʋ��,E�J#����W�Vlܸ��8/����K����?'����O�#0]�t��j�06m\�1�Sp�h�xA��1�������V�^�:�K���.�۩�

@f�u`��jąR\��OΜ����u-�hƒPmm-26��L>�DrsfN���������8���+IHF�}׮����<wA�e�z{�Ż644	I������^��r�`7n4z��I�P�� �P��o�-v�؉��z1����
h���0�k&�cI���j<ڃ�.��3�q۟��_�|��Wg��!���懱������׭_8�a����_���?Ѱ,��;[�����h��"9������K�M��o�1P�cJ[#�"a�%vL�K74���p��E�����$ڼ�m���/©+N���ޙt��XS���pR���%�����Уq���@��W�p]t�,doO�Ϝ�ɓ���عS&�!&���-��ၜӶm;� �'mo�@���4"f��X�V��Y����܈�Gze̓�P!����NMMLj��tRZ��餌� }ƌn�l߾ﾻg�q6.��J�zm�����8�Ν#�7��^���z-O[;�E���?���}۷o�@�6�e ���CR�eҒؐ>ٸ�\z��Xy��(�8|�(�X���c�Wc(U¯��w��1bHel�19B2ѿ�'�~�ǟ}�s'4���ޞ��_�uφ��[��u�OJ
��J�,�щ�}�Sx����W1�����-��.���5����L&�
!������[ZZ�¥P
--�^h���P�X	�ɸ����3���%<������9s����^���R��B�K�ƼՋK�Ago<}�D�% ��b�Ħ-�����H#���,��=o!sVw<̣��������)��a�"��B<���F����ILL�('��cb%3Dt}rf�!�J�)rRQQ�̌Uz-�DD�}���/{/\���h.U�d�rh����<���nkk�����/>^�����J����s�D>JJ���ko���F1�}�,�	�����Y�2Q�ufv^��Q12�^x��s�΄����I!��g�䄊�B���K�����7j��oAxx$FF'Q]ׄ��Zħ�!u�*TԷ�7?AAE+-]a��	wL�t"�������yY����<�ɧ����#k��I+�ԡ_Y����1���Af\���o�
Sc�n� �H�����YZYa�lFsG�]�%�J�����d�(�6`M�j������F64h҃�����#F�D�u��1StD��P�x&�}�J��hh�q�F>6���*DG� 3+KU]W+��|�R���Ɣ��$��Dn#K������z}�_��U����ފ��j����s���Fn���.hjjVe�����Ҵ�����)X(p���N�hB�aQ��mĐiTy��k�C}}-����	��J���٦P�pNw�wU��v}V�%%%��w�����ަ3$Յ��Q��^{��92����wKIO��������;zP^Y���N�߲i���������¼���\��o97�$���_���z��<�����9��h��շ˳��CNb$���o����CZb"���<;�)�n
�*&���2j���֬�l�
�qL�o��f8�;cz�ފ�cF˃9
���1�S�u<Ē�by5V:
K+��%�A� '4��U�V���O�l�����O�4Jug��{��&��jj���o��F$�H�j~nA�͖
{�mc����H�����Qsc-��twSh�B����S��������`��<�024 7Wx{Rsu	�~��56�`rr�v����O>�XƐ�*gϟQ#��ތ����n�l�g�ux��uIk���eX4>&�|���_��Ձ��,�B�]��[�����bϜ;��y3n��0�Z�7xu퓘�r�� F�Z��g���~��u�Le��x�����us����ъV;
�������<��#64H`��"��k��"��-�%�Cɠ�I3||�������_��H E����u�q�YaW�V�G#a�����X�f��B�������cH���S����ũ���ގ�^+��Z���R��s�x��ShXʵ�����^��8���&9�ބ7>6.Z�sUe9RҒ���Pq�x��!-)E�Alx����z�ċ�����B8��r����N��%�P�ڣ�1	� �G^Vu]�.�m�݆s�O�7^ŭ�ތ�o�V�����չ�������N��|��q���۷O�/1�=���3J���쟞� �*
��u~W\y���Ҋ��&���c��ݰ��{�.���]E�w���>���
OUD���7^.�n�0�l-z*�8�ؾ.߻� ^���h�*GBd8}}/PnG@�?`����ƶv�xxb�<_?���*̕�2`�>d2I�wf��{���a����ĲX�������a1��5�����nkc��ή.���8qB�h'W_+��/����\�?�#2#�'Ҏ����� �^�dT�frj֖�v�02jR���\~��d��IMMEdL��2%�2�!�VWS��0+3�M����
�������F`yy�>��vx}����\wõ�����(<r�&'�e͐Nb:�|�Tί��
���?��;��xv�.P�����Gﾋ5�W���#�j��HM�F[Kf��q��rw�Ǐ1<��P�>�9g̎ �g�/����'����?�x���i��²��u,O�ే���WhO��D !*B�$}qښ9]�� GF��Iqeh!�Hj/E�֯_����-̋��ǜ���U�����~BW�����`_�Ƭ�������g�oº��e$
_~�U\����ގ!6П��@,_cjr�^^�:��1L[�f�+JE�KL�CNN��pxdP-!�&fV�ͽ��1��k�76��t����}�#W���ũ����vRZ*��Q��7W/�|2^	O6�e<w�rsW#7wN�<�j������c��m��a�4����s1X�̳�ax���Q*B"��W��3�-:��C]S3�lށ�W_���4Їޞvy�m�����W���+���S�_���$����y�����ȉ����7������t����k3����܂���VW!+%~^������PvN�8y��t�풅�Y\����ض�V1���jy22y��8��0H$����"8肊���'�y�M�33hhh����1���2���D?V�4l~�E4l2��w�o���c�����d�֤_���n���nh��6�#�<������C��GV�*M�����#2/b8b!@��7'�Y4�ՋV̋�;Ї��Aц8���V�LΙ�U�T��ɟw��q]V����"���)&~����%�*�BB(w�q����7���I'����Ly��>��>�k�����޽����2ѮY�L�q�~��W���/��u�����3�<���։�O���7�j[��-s$k3�x�gw�ay����	�+��R0�ע�����Z��74
w_��(�L������+U�[V`�6�f�"=nV���ب$��*4,6���R���|(z���H����Ao�PnX���h�m�`�**���h�ԩ���r1�fx�322r�'�cغu���а	��~�Y��ަ�457���Q�i��uP����SF�<��?_����_�G����W�m�U~�)�4�5kV��O�"11N�;?3�cY�������x�8~����y�����g���r��Y����������^�xx���^��<�����ۃ�C��Ԟ�{����/>h2��3�}�Z�dd�o�±�����@T����>��m� ����W��-�|�W_.���>����A�9�����g/`uZ<�	�17gVn��ggW���� �2BLd�-E�ɞ����:cc#�V�62,z�I���Ј�t&��-�2C;~CÃ�H|-z���~����T=������N-S^A�6�������kd|U�uW�(�bϒ�M��V<X�"ٴy#:�;p��Y�τ�4�X;���S\�-[6)�^8����� UUpuq��#�gϞGum֮˃��;L������Ȳ����**�%�rTVT�7bDeؽ{�Ό�)��(���{��wߍ��6*�����epdHn �y�����܉1==���r�	�DIA�]>;�9��\p��Gk����{�)"��z�Ƿ|+))���_}mX�˻��~��WN�l�_���� ��z��������6�N�T賴X���0�`c� [;{�uucdrsǶ��!���[�!0�O�Ź�e�%����..Y�
.��^�
�Ř����
C��4�97'�����Mh�,�)���7�Th۱c�0*�J�B��ID�D���5u�YZ���7��k��mbcc��ҳ1�fu��RSC��G����ș�$de�[Ц�����$>^^��o���"�c���ҒrQ�SR����Jy6��<<�����s��]����b�w��(�P�/OGFv���:Z�18%C�=Xll���J��3��=��fx�T싋�Ab|�"�ݩ�'��� fĶm۰:o#:Z�0:>���*�����nE|R2^x�$>��|�,����zG|������%�_x�S�ֲ?h������7��.�_�|�S�4ljoe'$����ZۉS���G�FG&*]rnn�l� J	F�3�X�sF�������]d�&���0_1��V��I8 �����N�|}�''�I���c��U⎕��`uvr�rP\\7QyH�������S6+�4tVi���J��C���X�j��de���$��8���Mbk11hok��a/O�GF���
�����h�������Gl��iŦ�y��4�t544ay�R�olL�t��"BQ�X���y[N��S��F��D޺�����%l���R���'23ӵۨ�\>^~��XX��� ��s�������d��s���5�^��
���Sp���������	���hX�eu�O����O�:��׹iɸ��o����=����HW~�47'[{i	8��`��u--R�[���a�\�+f�+=#U��yl\	&>���� U6h����5L@#���S3u͚��d7���NU@p�@��.�;`���
��~��+:*}�T���]����C�<o%�oek�U��1=����N�Olذnn.ʟ�ڄ�;66���M�0q�qwv��ܹ3��O��*G��^쭵��X@�@�B�yb[,���B������4+OsŇF��ٮA���Hc�X�ӬF?��cl޴�ٹx��wa�U�;�H�g�nTT�!5%I�pa	�W=�}�գ��c���r9�b�K�̔�}�'��Xaإ�
AYY�(P�7XX���f
>෿{���C����;��↾ѰNU�G<�����Ͽ�j��?��[HO��o~q�և�ƅ�#�aGk[XP@��C�sh�hWÖ��ia�6� ^�����ޮ����e�Ɵ9#���a>�6�aa���QC"�<���[��2��0?�<�:����$FDcc���+V�HNID�_8Ξ��z�������V���eJN׮�ASs3j�09ŉhkxz�����U(nV]U��tLL�B���r�6YT8�yK|���i�)�qS]M �.�NF��Cؙ���4"��3\1�rw���بZST.��--.���J�Pjz���#c�r��FeE� ��n�1Qb�::p��cv��%�f^�������)�UV��Hb���h�px��q���r2�شe�<)/F���:;��DVN:�|�=�~t׷o�vjj��7VAE}����;���禦���CѩSx��W����,9X�c�d�205���n}@2�<��T�tJZz���p�cE���!zƸ�f5�nۺ�<������L����088HK�<{X�a!AXE��13M�ppr��=[P�P�sg�0=5��B����`||ˋ����CdTZ[)�1����خ���M���R��z(��t�3�yH[���L�(mD�d��6w�&��u��3�f����|44�)�f�oCYY�*�uyk%��"���[xSss�*Wj�3g=~�$~xFW�    IDAT�=ʛ��y�s��b׮���<aool��a�H��W.���>'\����kQ`:�Ĕ$t����w�Fu��k�*ޱk���Ҳ
�9�����߄��:|���o�ᚻ���s�UX��������Ϗe�$$�����=� �F����yq�YQU�z�RlЖ�~�������&WpŕW�`�i���'̪�X�WF6%�NF����ё!DE�&�ޯʆM�Ӡ����v�ns3ӘGsS�&�3W�����.`jr7\��|���?{Y9�����r��u!<"X!L���l9|���j���}�����΂bhhPF�m�feYy����s ����D�3�����N��L��Ќ�{\��N�/<,D!����Ξ���<|��$�K��_`�J~�b���| �Q�K�[|��n�e��2� nF�ܡ��'��⩐��?^R������\����>����Ȉ�1fd�p�\�����Ÿ����g{��w^�|���C����*�PV�����C�g���;��'~�����r��ҼT��Yl-m`C�eg�ڶN�&�S>���D�P�A�X�a�p)~8��ı��z z2�ff��;:8Ї�W쓞B[sff��P�_���#c#b�rp���)��DYu%�-�����~�D'qg(rqv�7ތʊ:t��b�b7�x�ͣ(/)������^�������#g��ϧ�z�_=��]��U�Sb�(Ǻ�fU�q_-Vg���N�=1�А@tv�ctlX�0@]]�[��慭[v���M�x�GƐ�6���X%����@��8rTޛ��vK/ગ��EY%�X���*���oN�jU����Rh�,�|�|��ւ�����L<���F�<�i2/�ةSg�c�n�o����9�i?�l(,���}��?�q����'�-JΟ�o�����p�
[+n�\������x�cS�h3a�,��%D�DX�&W�� �9ˊ�骷W�E�&'j2�����P��J]eƌ��0!�t���2Μ�\��Gp�w �v�P�`m+�#�&8���VYu��������WN�>�ə��~FeY!�|<U0�L�
E�Ѻ#�F�H�>"2�+��V�'� =#�C}R�����������_`&1'�'^oo��9arju5���ԐnAA�<��_""cT����#:.V���"A@�/*�K�������|��ԧ����ٴ7$%-!��%��O>�۶�s���IxeݦX��ŋ/��Ç�ܯ��2<xc_�)�I�ﳣ_ 6!��֭�N�y�����yyy#�豪���~q��ouuu�<��/�'���Z��ɒ<Qv��k[���6�����{lL�p�.�=Û�s�n��K4s+Q���_bQ,�	����_��\_O��f�g�V�pH���<<<�q@�b���:��� 45����K4;[%�darB��Rw����;gAaek����,� '+S-�O?=���-X�nŃ����x���ccCjwq��^���S%o���8�=00���lUT�q�UvV||<QW[���͛6���Z�+<2�1q� ��7 /���>�^��Q4��|<=ĳ��!Nu錸����K�;1>~��M�E��O»ﾋ��=K���lAm۾U
������Ι��mߺC��pjfU�5:��|�Ns�@�O'�������fê��z�G߲��ȹ妛��}?���%�c�a����Yႇ�I^n> �>JM���J?_%�4*Vz�
���vZ���vL��o�C�bQeJ�twu��؎��HJJ@O�1X@Dzժ�zH�-��6'��ͮ}Ww�򺤔dx��(w��g#���G?="Ȃe�<� �t2zU�M��Iu���l(��P���.񵄄x{UUr�0�9��< Ʌ���� #1���P�$�G؅�Vsc�����p#V���Zm� ��ʺ��Tjun.F�F4�A�%z$
�0���tv��ǰ:7O�Ӡ�_���O�����x)B�,�,�yQ���P��gGT�S��C'�n�
��E�e8$i0.!Y�#��M�����t���?&FG�_y���}���Z���G:ȣ��2Ӓ���,����s�6O����1y�q�A�r���(�.�_q��h�t|B� �g�Bf&�����Dz�qS�W�E��/�/���D41!Y���CV�+q:X���9U���M�kh�!#5$( �M���r�k�N��u3��;:9�LLHR��y��Nxyy�3�p@�};�"O/7y*bT�^���H�������_�R}�G�g0)���P���\���Ubp���!1)M�â���!;'����7cvnʘ(��R��OP��9I��8��H��eJ�7��2�8a1��s0=ׅ�jk}��g�2���Y$1�!7��#�?������j�ؗ'T��ݵsgSrR�.{{����[���n�TUU�<��G_ٶm���&����X��7,LO�Z��H?�F�Ʉ��E8�{���������AÑN�ܜ�t�t�����ʪr�n���#��%���|0'O���XhX�$���5�<19���PlشU�U2`np��`eYSY!�۶����#4t�&(Bjoq_ǯ1����6�*����`��"-..DcS�4N��W��y ��	��YX�(�ڢ�҈�w�g��"���+ݫ��RQWXuI����X��
�N�8u��:�����bb|R ���� ��yy�#h�lW�Ix�a���)az���w�C���E8�b�*]��c��y��b�p/6���1��|���?qJ�mjiE\||��7:::v]ְ***��~�/�����_zE�v�*8X��qXrۻ���m����jpb����߈�EP����1�oL�d����v�>���Nxx�*#6}*;��|��D�痱e�vi4���KX�z&g'��R����ڡ�`�916���x�Y��҂"!�Y٩J�	Q�:s�7mEZF&�q��IDG����S��@hcc- �a�?yb6V������bb�����)~ӎ�[������Y�Q���Jy���7J#���H!��T
m��u`��������qM��%(B��8��X,c�0'��c�y)���*tjC���rp��?0H�v�4ll˘�����!�B(��WTP��_~Y�yN����;��|y�l���2R.]��m����]wYê����ٿ�}Ǯ����C�%&���bs��\\�{��%Yh��G���R�040�\��+�4v�P���5~h
���Ò���"����)������k��ZD=����fM��4�;N������݅cǏ`|bN�N�b��0O.���NOᖛ�G{SN;['Q}�2���R�ƆV1��h�<g�h 99�u��81�۲u��l�o0�Z�v�>�]�}������a\�p�\�����L��2.=���x���DANz���P�ڽ55�������-�Ӓ`�@ͭ^C�"!�E�������������/u$���?b��+�n`��Ϥg��]n�$�����0��j�މ����s�������><��38��g����(�>q�
)N�[ZZ��رc����۰<����c"co{������ђkp�a��"�-�uga���.�&F�OЅ�(����xx�i`�v�t��Ri�P��y��W�c�,����m����,��	���܀�ɑ�ʊb�����U�s��(����4�7!%)M�aGW�0�͛��' ���]�j04j|�P9H��MMM�1�W��uk�"8$�!z�-͍
���45��j�PN����'��¾}���ت�B��+�3g�ا���rD�#UiXA!�8�[�R�[��;"ʐ����؈�{��e�#�3/"�[|�$D�@X�ѰB�#��;�H�I;�,�Uʯ��/�+������_�R�dEE���kfffd�����GGn� Ҋ�
���҇&���=����==\a�e�s󰳴�ȄG�؛���D8�[�v��E,������bb�
�����᭢c������3Vc�3.��u~�/��,WM��;+�,�oh1��B��;��b�
���w���8�8b�ޫPPR&��޽���~9yM�
Ë��=��Tb|l
k�6H����M�>.;�
�I�J{�ǑT�ih�l쇒���ֶN��#)!�܋��B�T�"48��	2��V�z�M�Z����#vn�W<٫r�/�U�����Da����_ɒ���~%Ʉ����������OL7����ܬ,�]�r�w�|/���"��~�3!�M*��������طg�S�b�__'�'N���5��8�ũg_{�۴�T��ZaynZ[����5jei�љY4��ch|!��:���£a\���2�,쿆h�L��&��6�U"C��փ�{�67��T�М���s�v45�kގyBvV:F�{P\t�n\�{XX�cj�|�����w �b����������Ҳj�"{�*��y(����׍%��GLę���0K[LO�#(0�	ih�hFUm	�]l���%����W���iz��X��
Y=�Z�	;KL�����
!A�HMJ�`� Ξ����(U��!(()���7���11=���a\��#&���c�E
ϕgJ��%s+A
�˂d.E^�����T� EhY�������g�v�9���{Ժ�4 ���_QU	�W�������������#Gnx���^���g��k�5�M��%���Z���7:��	�c�HMC_o�n
×�@++�QL��%y+> �"9A,�tZBzO�vl�£��D'���ˋ8�N��LNsWe����:q�9���0W���˨�b�ηp�d����Ľ���}�������!�I�����#g���@��W"P[TX,�@_� 5�	�.,��?�#c}������P���!VN���Rȗ"��jI�E��2���T�����c]�z��V`dpNnؽ�
TU֪��
��������"a���FlZ��q6���i������f_Q�D:{�@/_��'&e�����A@g@�RDd�H��>�,���q�=?���Ey�y���e��s|����wDEE}3@����W��O���P���ٔ��*^+�p(�
]}����|)s����Lf��e��[�7KCo�����[���o���m��~^0�r=G Ɔ��kٙYHN�GA�y1W�=��X��ioQ���%�8���73;�^����^w#�����
++��݀����6�"�HK�"tsc�g&01>�x�+���k��c��r���Լ�P!!~HM���� jj���Pgx/*(AhH���}�C8s����i�S3�(�(���=��\aog�ٙE���?�b���WU����)iZ�YXV$(cǮ�}s�aBl��ҝ=}�kegr�(_����D�T��6�*��k�P��0��/<��5�\c, ���gt�n��v�ڻG��9с�f����mc��X}����?��+Ã�α�Ѱ��Ԋr�����-.[����Ұ"���١P�C����Qj��=? C�[;�vİ�`[i���a��=�7�������?x�gf�Zm��l����������#�cb�9p��Y�Lϋ�@����a��?g訏����5��F|\*6m�%o��ӊ�zU�ӓf�<��}ܱo�^u��K�jd�ujH�`av��~��Z��H&��5�HO�u$}�2�#>!I��h�oS�F��hko������uy�-M�Q�nڸ�����F������휜���韛hݝ]J��6����9�]X����dm�%k�g�aX6^�~5��?���|�%�Er L�9Q�v�F���Ȱx񹈀ޜv�駟J6������/���ƛӢ�������߿��;~���^�Ĳs��P�dr�6��kv~Y2�����S�Ƕ
=8~ �j�d�	�F"��B��&���1�d���~���=��ۄ:heL/�P���*�$�j��\-��n������3�fRv[�[V���|������td���yb�U2a��՘��4�e#��Ī��˕�{Pp(J��099��k7"""
U���EZj�0*��L�`��XY�FQq%f�V$$����X-���Y-2���#zJWg����ظx%Ԥ s��$�h8/@f*ϔ�s3�X�R�Ғ/�T�Ֆ����E��w�vR��Mt���𧇌�Ass��o߱CFM��=W\)��s����Zj��56��֝߾muZZ�e�7�8��x������e�%щ�O�I�u�g��Ձ	���D���Ӈ�n�d���5�����d�����ݻw����g4�05e�C���M���N+=��SJ��C�EF�<5/(='�q>���RlڼA�S3<�{w/�[�	�N�Q-.:nھ�j�LʈP����Ԃ����Ǉ�[)��n�:Cnk��̴�#��H�IH���1-W�����0� 3+Ed<�҆���������2��2�`�C˓���F�l+� $,X^Z.e�{��p����b;q⸚�T�fo�?�H?��P�Isr�hX4��'��y����\�́��{�1�l�!��Es2��&��|A�;n�����W7^ְ^���z����]�ÂB��8'��	)�q[����S�pvw����Ձ�`�;шHd�~i;֥Ig�bX�����7v����#F<�ȧ�F�x��AyI-����c�@%�<z��+�S�l��wv
͍����j*��qEN��ٳ��'%$�������9��$�%����#)%M8�[����$�^����⬬x�ڣ��	����M;1a������@BR"�Z����K��WI��b�)I/����`��5��^��|K����j�A��WG����[�������(}|���)	���{='`��3����'��ɨ&/U䛷l���7^}�%�m۹KR�4xVצ�y��������.kX/���Տ>���ޞv��Č��x�V��ə���2���9-Ub���ӭ[Ŝ��+?�/���C�!������]�	�o���ja��KRzZ�����U��S���ډ��>��8
��h���3��͈M�Қ�ҲB��7bߞʍ�Z[��щ � y[rȘ�s�J�s�a�C[s5b�������7#=#[=<����W*�\�n�YbS�(�qQ�1j�rK� ���`tt5u��-��upv@wO���{�v�b	GdH=�e".&	Ǐ�VȻ�넁Q��à��K��&P�F3^�m�w��/�c�-jIQ��0�g����s!���C�QL���䈪F�0��3�{6m�O����׿��Uk�p��7��r��4,m����;�]q�-�(���9�����{��W�"�lm�cq�@)�88`�<���ŭ�̏��e�a�zIu��O#b��8�vj1��f�AWG�ʳeg�j<��~;{[\s�D.ZZڑ��
#���JJ\r�@WO����z�We��W$��s�A��* ���PVV��z���#��X�[_�++[�Bã���3�%����->s7�7nܠ�A6���ڰ~#lm�Q������Ρ��A�n�C\YY������Qd�f(�jl��4x||,��b���&p���	{��-�E�����BE�剄SI���N���F}}�1
g�M����9�!��5�?��c1#����m:>K�B����!���}�{�vJ��GeXJ�o޵��}�7��~�� )���z��y�Ԕ$[�͸9;H#��aQ(������3�ʱ�I����-�$zϼ��vfjZU!�X�Q��� .!F�:Xj�����a���锇�1��TVV�yL����`dԌ�%��w�y+:��q��g�X���=����Ț�����9�2��\/՘5�9��rAyI)疱v�F��y�����i�'�  4X��5�u��	��~��s�'ùr�<>+�q�YRǔ:gϞ�����.8�Ҿ���DE������on��ݻTᵶ5i�Rvv&|�=��ڤA[6��	x�r�*��Mt�}�    IDATb�[��I@���M���_:0$H!�8!�� Q@��6w3�y�����Px	��߹��4�Pp�<~���!0$TC4,�ã��Zp���];�ڹ9����瞻�����Z\L�=�����b!|�T��B�i@��P�^� A;� Y�%0T����K�;	�쌥�ƶ	~Q��"�o�������Å�|���	�lmk������r.{;g�Whobb,||=��X���J�'�a���hjl����d�����0!�C������������3ib9����%-�����(����qNt/`���Ԛ�[����b�r diyN}���q��Vi�#C�����0a��yV�6��@{�тr��Þ�;QTxA�CN���M���|�hi�c�X��RkK�e�U8t��E�c��˽XDM˰8�!��2�:'����ɿ�3��Sض}�
2>�>�(�"�T0�@�vYi�ٵk��ܽ{K�e녿�p�W=�FDX����;�f�m_�P���6=V�`��j&��~�Ӱh0�r,=+e�yCX�ѨX�34u��������
o�{&���U�)�-g�4l�U�p����k)�6_/w���T�{y�k����a��y�A���#�
��wȫ�#P!f�νpqrAW5��T9�����/ �DĶ�V-�U����y�J5Cz8��ҥ2Mtt�������	q	���vk�j[���/�������HKM�����VS��ø�Y���b_
�wVN�6���Iqn����k	s��FFFhW�T,,�(��is�W_~M���=�nz=�X4,z�'�|Rw�"�@�%�wV���sy�6�up��ˇ�_|��G~�B�|�051*q2���m�mnI�5:f�+���j���(��k�"`����s�v\������k�������n�I�U�55���Y�F7�1�E��s��'�=�����+噹�		�qq���k���X�ё��	Ji��)��������N�Nѧ�\��Cf�A#��a�<cc��y�:��cc�<����iJP����~^���Wc�#_�p!Ar��SK��r@��V��i�|jJ
��XnڰQ�O�C�)���k��9�ឞ^2���c��lx���K�^���朤/��YZ*���/wOTCj�%âX�a����O=���(����PH�b(<���֭;��w���W���������\��11:$��-��8�D��aXn^�2�֎vU@(i<��@�Ke�dh
b�5l.SZ�O~��,��)$�'a��]Agxsr���������	�����PK��z��i�������t���4��βn�z��ŕ%���RR�����.���
�~��'����k���KPvN*��!!p#/��s�X�����3Z��1>6�M���QZ�		��T$DM�z,,-���_������U,1�!m���na�D�#҉��Hg�^�E,���C��\~I�.C'�-<<ܵϚ8�-F���}/'��,>|�#�b�/�BF�K�Eh���GbJ*~��*j0�'�Ei�3��v�����{��]6�����v��w�����IÚ6�iI�����7���@o������^Y=-�o�o�I�/~ ~у�[1Y������1#����t�6o�(�z��� Unu�Հ咠WWO�ϭ���Ganf�7�W]��$��֭�5��^��#��jM��N���g�hia����>] ���E5t�
��֪=!%A�`�<3LS������j5?sp��ǎi(#!>s��(-)ן��6��R�}@iDRRRR3qFXP?�#��h���J����"ۂg����Ks�|������)B����3�������ó��QX	�w0�gضU�s`�F��=?4��gω�VZV��e(��а�(��PH�������A��)��[��_�(;p��߻r����֡C�6�{��︹8��`qnZ����P9����2,V�܄���B#�fK�1�=��� �O�HY�0�OMO(tw�Ԁ����V7�0�$���ǎ.q���xxyr��V6Zm��T_/��4��}�i�2�Ƚڽ{��i��7ܨ���O�.�D��ǀ�摖��q���"�vvsU��$߬E�S�R�b��̦VCdx0���no����T0��PYU���p��,YXK[��J]L�ɨY��AR^�4���y������}�fm{�`�̜lKL��rC8�ȑ���͖�+W���	���f $$��#�ّ��rx�ω�_�ޝ�%�[/�ҹ�;�|)�Io������Jo����۹�䲆u��������--������a�e%�L��VD�����������d�1��r"�އy��F�A�+N���W]q=:;zQ]A�aW��))��J���SŃjj�@sS�b~vv:JK���7�o��^()-:L�ӑ�A�'�$^FH�m���5X�GDG	S���u�e>)�t�\��*7G:���s!�)�̅����"ͫ��$y5�@���dgWg�`y��-=����9LLOa����,�χ��5r2���g��݁�[��9w�X�bL��`���\\UAK�/�{���O�:�_<�������h/o�vP��kw�Lf�eg����>׳�Pp^���׆������x�7pӭ�	y����YY�*����r��޵e��R֣�|���!���PX[{b�n�zY;M���h�&&'�53 ݂a�R($�"Q�ZFG���b��$��Ŋ=:�{��6oވ�@���DH�OHH�����AHx��T���ΟDX8���u��nW��z�8q�344V���]U���8v
�6HNɐ8~�(9	�Qpq���S����Wgxz����VJ1����5������Q��i�䏨q������f�t���?�ѱ��m@kW"c"����A�nMI�y�8ȽgۋMu�N���楼��UU̥.==�8i��%����5��L���lc�φ��$Ur�:C!����!io�ubXhX���>>_돽�ꫢ�|���`��2f�S����܊���7�~�y��=��XG����'�~����'9>Qp���e��C+��;�g=LF�&��*�c�1I͗�w'b�e�EA��\��	��Л?v�B�-�ܬ�UVV�.}tT�ɜ:�m3�>4�5^�����x8�Hw'���-p�ȗ 8t��7`��M��jo@TT\�e�]�XX�@pX,&��Z�9aGX�?�<051��s'q�5TU�����ظy�F�斖.2�1�W��`��tOO =8�K��t�����>pquWA069�؄HU��%g����Z#�FQa�
j��t����]�'�6�*Ӊ��h�E����L�=����hli��G��f�Fϳl���A<FN8�ϴ���Q9/�O y�Lk8s���^x^ľ��k׮��<s�f��05���-7^sCHH�!�u��!�~���|���Ǿ�N��W(d0�Ǣ1�_+�YXBOo?���eº��ζvVH�!uM�X�0�Bz�!	e%��ܵ�ҕ��Ğ�*�
�p;k;|��ocr|R\!�ҵk��߱!���;;��y)T46w`�<���dD�����}�m�L���UZ ��Ճа8�Z��O]@o��RR%�A^VWW�c#`cm/7�wv����vNHHJGcKںzE�c5�Q�q�����0�Jl���>1)�vN�(��DOo'�g�1�h��X���|�|��; <������2xD�KJ���� x�+*�u��xd�2T����)zb�`tv33�_N�L�6������B9/���<�}|͸�8������5���.s?�$�8�����.��m���۳�/kX������o���K>$�9;�J���ɮ�XZ���Ҋ��IMRrKQ|�G�����;?<o�%>~�ֶv}�D��&Ym��Q����Up �~���L���	cb3)�����
Í;{b��]hhhAQ�x�8!5)S�Ø�����(��������Pܔ�ON����
�}�X�.W"҇�[�֭;����:�u�����.�J���s����,m�(��|��z���KKK���0�M=��uENN�<PO��V�Qm��.��������0�`��X#�%����	������"���6�6z8yμ��q���C����7����)�%�aP��W�'�د~��<����;rWP}}#��Q\Z�~�?6�[�_�������{��_~��'|�����+�i���I�]����jw� Lc#pqs����Y���F����p��p	��ЅyR����a�	��bI��썙'���B�f���:�.joG\|���"mĺXJ��'!19���?Tp�ڹ]���M�ڀ������$4�u��4� 5s�����%��`��1!V~�^~��FQa9�m���)n�-U��ؼa��QVV���ARzU6�9������J�,��Օ�{UYTu8a��;ב8�ss
mG_���/�\L�I'������������&p,�x_�aS�~������XH]Z��ѺI~^oo��a�K��#����u�]*Њ�˴�������g��뮹�A�.
_���7�99���}?�sqt�����}>�5hX�mXZY��iT:��{�@�\D��@�F��_|H�Ľ8���P?s�� c�ǻҒS�Y tvvi�0,,\�7�%�w�bdӚ	��,�'�ٌ�� &7�!4$(������yvVTe~���$�{�p�UWbj��FeNz՜�VVv��$���:=/���"��{5�H��Ξ!ɑ�x9ٙB��{t	�������:~�		ؼc/��eؒ�����h��P�;iP4J��qE��1--ZhX�|�C�)�4�HV�N��1��Į|t��w�X�x�!Rf��E�2w��T<��s�\�����II7�h��[��έ[7�yY�w�c�~��iII�?��#����=�$���0/�"�K�kbrZ3fܳ���P&�A�t���՜��a�|I�#)9E��?c.������o?�L��W%^�؈����y�9��F����I)\Nl�Kyp߽���-((�@�={E��X:+�]۶�����
�+8��1+�6�#�wi�@4�1�q�6m�����$'�(��h-	{驢ɴ�5���n.��ҢX�d�z����; �}�46/�P�xaNoCڴ���E��H���͛����ji[P˝Mv���^	��5ɀզ��eC���Sސi>������l�)_�tӳx睷�{�9����c�)�LclΛw��smfZҗ��+\YY����?�ezr�/}��uEy9b"�&T�!"fi�eJsKKZ���ӧ<�^�����ݭ$�7�����h�47��$��d̷�[jcm ���q.q��Q
�/�0�I�i�hzLT4��je�������,"©����%j�b|�M���_��Q{~���
��b��eK����Phkkm�`723R�+�?����ƤyF9���DI����	1ѡ��1f���p��㘚_��E���Zc6@4j�(�����E��j�����N�ǵ�7��^��k���\���%�=*ϔ��gȞ�y5յB���X	��f���1ml]�~�����E�RW�L<p��v/Κ�cbb���W�+++�����"��~���l���_C&�ziD�Z.D����	`B�������>0`&�+�fX^�Z��0|@�8�b<�%�+������ػ{/֭[���z�kҙ4#,�p��U�{�#9!Y!����g�e�Ftv�*	�����5I|�8�e�]�Q��\�m��M���D_{7�*����
�<5#9$k[[��䚏�`Fh�?��Ŭ%nE��ݓ��㨩�N�>�2\;gi�k�3�7i��-��АL�gQXZ
7O/���08D�/c����g2Iy���k�
P���C��{~�S	��`cnsڐ'�)XZ�����_�Ԍ
�@��K��Gj6�92P6�����i�W��%ģ��]�Gg�p�fb��=�N��$$$|��;���~���Y,�޸�h����QUx�E�h��jq�G�)i�@u���I�b�E�P��%0�E,�FE#��������;]�d�6
����Au�uuje����������R�}l;�9���h6�[%���$P��c4���.�g$���}��i�ERB2B��5w�����p+��\%I/&*�3(.:,�#*"Lr}S'&g���p��9�;���Xx�����ь���&�o��
���a�07/H�9��ł�H7�^捬�l���h�5�k�+Z�{i 4&-x���z��P2vn3���iaq���ܜ��� ad�we�98,D�kR�;w}��o=��ݹ{�BNv��ݝ-o&&&v\6y���U^^���o��������)$��hM�̔Yo��g���/�.�����N�>��δ]�pl�0����f��0�d����SE�[���x�U�u�l�f���NN�%�9"���F���S+���{�,�w�BR��]��]|�p�ԗ�La�aZ��œ#�����~ >ge��0��~8�� .&>ޞ�;��!26Q\s�
���8(w4>AB���u>4dP�����=&��"�'�m��&��e&��c$`�����ǭ���[u��*����	��i�4*�g,�����#ՙ9$w�P=�z�4,z::b�T/|���{�^c���N2O4���^�4�˓���hoo�7//���_��}��ǿ�����KQ�y|��ad��)�$��P�K�Q�c�nJ/RQQU.D�����h��>X�r������A����k�����[�a貙3�ְ�<s�rv�i�U5@������Z2O�r�����6���a�����}���HCTD�d��:	�)HLN����0wkiiFKs�<8!nf��X���8�#c���vqM����j=4��Q�΂��;��Ƨ
��L��t$G�x>��4���B���c9�C��qx�}X4�@�ת�9*����V$��_�0J'llWpe��eoO�v^t����`9�z��	�q��YS33���Ru�/,��䬄H�F�Z��Z���=G.뱞y�;~����x�w�x����y	1Ѱ�������L^44E]�ܰKLLM���\�I;�<��n�A?�0]�1PY�C�m���0��m[���� *��-�ʑ7����w���q�6z7޴۷JV���J��l�>zT:�yY�hmnąsg�� XY.���#�6�T%&�����E���_��r:�ʎ��y�X�
�f�*?�/�;;���\�����r*���4iȄ�I�i�f��A��#&����hnl��j|l����)����T��a��U,�3b����X5�����-[7�(�l��3���/7[5,>��C�+���czj��:z���@Ҝ���2��o��54����.��� 08D4��¾�޾{n��w.kX�}�������
v���ƃ�'[[x��薲�X�[�'�a���8{0)�,��TΝs7M�3"�(JVA�0���������������u�Qg�UTL��b@ń�HMwӉΩr��;w=MɈ�w}��%�T=�<���O��s��"QM� fa+���w��Zx(��s���/w+�4�ܬR��SrVd�I8��ذa�J����Z%�,rjT�P���Ϫا���;���W'eA�E]b���?��s��Q9h�>xP��-���'�Y�~�,X�H�>��ڽ_���g�Ҡ���_ʎ/����l�_Ƶ�"19z�V�5��V�:/�7-M�
g�'4��p�I���nڱ�q��͗���n��@̈C�݈��G����M,��U��5�k���j���f}��gN5`2��T�s _[�Nׇú~����š���O���Q�G*_�`��oi�*M�{��Y���믽Ҙ���Z����N	����˒??�����T������jٵ�̅�ъ(SU���Bz�!�g�-�D��*3eDN��?X��T�����v<B�ǃp4�2�    IDAT��g�ƌ�ׂP�	��-^|��w�a�HT큒�|���[�d��j����[*IK�eP�`�`?v��h��[�J1��"��e7��AUP���83�%�fƌ��ߞ��>�_Ǝ�(ë�+h���+CG����Ƹh��O�3��t�Cw����R*�Tj+G*�	���p����R;�QQ��b�x������2��lٹ{�:-H�M￫��ر�+�Ե�*s�M�`�,V��C>�c�!C
h���9��tV�n��<�`C����ސ��ٹ{���5�mw|G��ˊ�O-+.��u�-~����}�]�l����������;�z�Q)/.����BR��k�-�@([āwH�F=�ťf�;�lX8mDF=b
Y�G��������D���fj���/�T�lۢ�� (���jV�M��v�Q�j���H���m��њ:ٲm�J��G�7���'�-��+�u��|�^οp��rK���Y#ݥ%嚲����Cd��3��X��R�֩��y�(��~`RN>c��(��G�u�3 !�Q�FT����aLHT�+�uR�]���F*�]��:@b��� Y~��?�7o�����s�IWG� �B�^>��̞���]�+!�m�	~P�4=�5s����{�g���
U����=����7���R�������^V,}����g�u͒�^;%��������V<p {�E��K/�_���X^�~`q�~_HB9XI������|n5��<�'�^K��8q]��*�裀M����������N���d�K=��`�2স���Cn��v�	e�/���o����wɎ];�s���EM��֒���R�/(�76}���O�A8��4(���4��7��T#�HtcT�@��_+�EL�F� Z?�=7�P�I��4_F�������|�[�$H��T�h,��뽿�C6 �f��c{�ٳK�9�l@����� �z�v�@����O���?�p�s��q����'i���/w�8��#�\���� �����/�+_&����������M�\�����ߗ_��ҧ����ˎǢ�_�#�~�����2a�(�S>o���p\;�9\��5%^����������U��-Gd��	Qy���Sj�h�?�X�8�Ʒ�V���.q,N���W�46�����پu����x亨��,��"��Ig:*�Q��E���~6�K��s���B�u�S������q��W�<ҭ /G�Hs:���c��������$+ �\6�'"���m�a�O�f�.�W�M�����t���g���ix��;5�R�f53=ph��`?~����~���ɓO>��U\:H<�l9��	2y�H-�}����x[��0Ϛz�447��77HYq�Nwݵ�Z~�O?�!cF˃?.�mڼ������W_��)�u��W�}j��/��������JN;\~������C�����_:;{�sN���JVn�J��L�jy��� ��ۥ��K�3��֚�[��|��#�L� �9��/���d�mZ��L�B2���TV&�.�Tv�?(k׭S)�a��M��L��s����Ͱ���ɰ)���� a�x�9�D���TIEJ�(:����HI9\�:��E���ä��A�ؾE�c;�4���-M���իv#��ِ���\�M= oyy�L;w��_'5�����b��(�ۈD3���~Og��ɍo��a�i�o��G��*� zy���(��xJ�l�p�3g��|Im;��{�G��˯�Ire��4��u9�G���#��]�����'�?�U�n���n��N	�?���~~��������d�J��}O�z�!9VsX�"�hB+Db	�X<�Ã(��a�+�S��y�D�l�d�9��-Ǜu���;o��#�?j��������dsbtntC}:��S�����ԛa�����:ݜ���+vT�T�dD���I8��͛?P[b��!�z)e����x�t��HmM�0��y�ހ��{��qcFK~n�7�i����H_uf��\)E �5�Eȭ2��pu���(���=w�I�BRq�<��ݍ�h!/�ENi]���DJa[YE�H%԰�����D�c|��ꨜ6�L:�J��,}�Q��k����/�2z$=l�C���k��˭w|G�͞'k7n����@�9|�5W�|�ճ�?����'�X���u�h��S��w��-!����r���U�b��wH�^N5 M�}�445���B���Ԗ@j�JG�+]@�z�{v��@;kH!dʏH4l�P��$��&)z��y�w���Bf��Dx<>Ge��5<2(�B}�8&�����X��&_c7�zH�]!&����.bɨ�A�$\ow�JF6�z=BP`����d��~�i�ޑb}򩄲��.T#�^XR��'{�}���nBZaRl~�C��1cTC�9R��f�8dH<��[+V��k����ث��B�s���ʒ��G�����~�~�k���т�C��Ȳ'�p<&?����;�HY��·E?|õ�v��O�
�{d�E�V�Y][�T^u_�L3Ln��
�����ǥ�}�,���^5�.�����wu�)àD��>p��bhXox�
'k�	j�a#�
����nj2����ëaqh���jk�ʤ	5ZNc~�&�xG���4#=���ڮ� 2C5��ۥ,�d<���xr�_;��'.�=c/*�)+�5mz���њZ�M�`0�ic5������oL{%޷[�^$��0_�����5��r�����!��͟�k��+�����A�'B (AO�_^���}����r�d劧噧W�W^"���5����.u�}�a��+�o}G�m�D�xv�D�48��}�U�r땳N]Wx��+<���g�Z�lB"�/�u���o��W_xF*+*ts9���a4�Rn��F��2pQu�x��/���:���l-��P%�����3�A$�EeH7`�o��3&�92�)� TA\��raT��>4z�3 �Dl��fO>���Ch�{��qzm��hB�%������\UK8|'�Y�0���;N��ﰻx~���z��=*��8ޢ�5�f0|��'
 &	�����s�齟=����]����=�� ���|�r=Կ���5�⠣����MP� ���~���o��:9}�ir�X�|�m��k�4�����[P([�F6m��T�%>{������;��y�\!�zl��g��;�4B��R��P#W]z�̝>U�z�AID��(?W_+�.�����s�t��̢ v��P���}�YZ�k�2l6�����\��f��x-/ה*�+���R�-��4+�0�7���n��wޮ�$�$�~$�Yxzp-�*@ӱ`�w�������/0�s�H�vs����ڝN*���C�| ��9 ��0�f��C��#u ���6pϰ�C�5Ƴ3Y�*rz�����.֘�`�����[����A���J"�'�?�F{|�\r��r�-7*#b+A\��Ͳl�
Yr�Mr�o�u�~.�=���G���i�q��o��峷�:�����\�ܳ�[��T�8$&�v��'?�c��u/���R���f�n_$���7e��MMz������P���؆ @�1:27��kz�J* �J`�8�����2��5��J7����B��CGnik������C���x�R@L_vz��N=�LI����W�� %p*P��P��H�@m���B7�#�l
f�t����O��Gꚼ�8#�d4� ��W`B�v���%�/����v� j�y3t-�ǰM�`�EG�r�4K�`r=�����Xحعm�[���=$[�~)?���eA�ڣ�嶭R\T +�.ӂۻ~�/R>l����*yi�f�JL��pێ���뷯��������V-Z�|�3G�Z�v�i&������a�}�r���ʣ�Yzښ�% hP]�}}�?�O'c��)f�Y $���>}0ʥX`#\�	���SC��j�#�xE�q�㼟I��)���,�O~��y�۳W�ƍפ���t���s��k�F���j7bS�V����Ca#�D���D%���|�Mj�Ca3�Ν��*
7��x��\(�&GJ���!���Tx�֭Sﶼ�L�˰oR�����eݐT ���5�q��\��N ����x��T>w�p�NSݺ�K��{� ���P�e�&(˞|B���Z�f�m��ǻ�O��=5-2h�Dmz,]�v�pɜ�p��o �#+._��ŕu�Z}6�O�M��.�p���5�O~�IF��UKe԰!Z-B7�(�"qc0:�J,!�L�p%���� �H ��< ����,v xl��h�~�'���c�Ш%h6�?����WTh��\����ͣ�ߢq���5idB۲��?_#�RT���P#�`$U��1-�`)���3a���M�D�?��#9z�F�tt��O�)��{瞐P�	.3l|�nh��A�Pm�axc�B�/��P�XX���X�<H�!�h=�` 4�1��z�y|.;/O�RR��s�e��e�5�JWOT�o�!�W�/{B���������O[!Ͽ�Y<�%,(�X�Gl}ͻo�|�w-���)%֟Zv�ҧ_Z�����W�P8�1v�=�[Ι2Q�w�yf�����$�:��]��6��dJOdQI��W$�i�p�C��Ԑܺu��g�9U�dMc�-�Dܳ�V�&��}�Y0b94�3�B_������/�S�H]N��Ӧ����rO�0+��b\R8�H��w���:G�{İ!����ݥ�h(ϴ����מV�Bx2��暈@��A�P�m�o�n΢JO��\�m�����%fu��EG�B#���P
���A`���z	HP��8R��	�� ᯑ��@:�UVʄ�N�a�%��7��nYr�2d����&	��e��=
�[n�Q���6ٰi����O����/*�P@\���zv�p��[~�dީ������,z��c-����+�}/E��d�[��~�V=�B�^���^�ɧYE���b1�̉�3N��!b��>~�X=5~���g�y3�U%���_0X<T��-�CҒ�J��&�b#�F���Q�%��4�S���K�
�����k�r���7�=Z��Ŵ�K�!ZYw;$'�Ic��Ї��,H��@����D�y�ŒL�ڂ���&����cP($9����E�� ���:�L���J"İ(x:\%2�LP��F *Nv�>�yy�}��SQY��ֽ�a�D򃻾/�'M������/�e7m���w����m����U>��F\�RI�=RP�/^gL����o�t�?���T�ߖ/^��e��
�uШ7[B�����'�Y�"�?�@>|���h�+3m��͔z
$��G���A�c�(�=Z��K�b��ӕ�	0����M1 �#��<L����Q���Rs��j�p}�l��iW� �^�@�Lmln��3gi�!����VAt.�J���g�A�>���z3Νn<R�_**��j�P-.���ƖF��:i�Ʉ�Hu�za�J
�.<6��b�3Yv��󥱱Im*��I��>ߢ�9|��b�Ғg�b���d�vܣ�>�������$� � k^\V��T���,�X��Ѝ������d��?��Oe��)�����?+��v�+*��Cʋ$ng�}׍�͹��]�唪𯏬��U/��i�T�K#���R�>����x�\0���M�ɪeOJs�����ޥ L�L�5�,$eL��<��Q�8\��}�T]H�ˡ��_��܌��A�ۨBN��gL�ů9|X�C ��� 㶼�T��	G
VUUJ�y��h�ТU��S%S6�T\9D�J *�TU�|'����F��ʖd��!�*���Q���u�٪�yNT���ςT#�C׻��f�� �q=t谁�a%E�j����ʕ(ܡ�jj�FH�R�����bWaR�`=8��۔�6��w߭Z%ަ���_�R�@��˗�4����ʶ=G����|q������)V-T c%���^{�������>:%�|��EO�z�����8�bwy���IgW+cV%�LI���t�ʯ����]6Y��U�x]:%�����5�%����8�Yغ�G�$c�1Bk�ּ��ģ=�S&O����ba !����X��j
��u�@KS�*�����U�k�;��5���ϷnQ�S��i�d U*;��]����]&M:]�T;s�I�0���vf����1z�hٵc�N碷D �'ͭ����A��r�7C�x��!�:���3a{Dզ��}��� `2�5R*}�yN�����$��T�\l��yV�P9D�@0!�~T ������'v�GhŬ���ԖL�vT�>��Cړ�NɹE�r�o�"��~(�`�Dl>�C�����+!�����_9��_ѩ�Џ,}�G�=����)�r�لx~p�
�s$�u�ϖ�(|��K~��*;wl���xJڇIL2���'ݚ����xJ�����Po�t�S�����O4�3w�l�q��������?���k�0|n%�Hs�O�P&&�m�:0I�D1�����| ��揶({󒅗(���eC��G��w�R)���xR��Hv��	gd�h��F-xE2�����v}v ��@��TRPUAQ��ܽk�^��16�3	�^�g�`�q2^�����Ŧ��������� 1�C�2ٞ��!>���Â^\f�F�P�@C|��vG�9g����{����4�9D�J%j3�h[*!%Y��NE%�w���Wξ��Kn:��zdٳ�Y��s��6�RΠ���$�j*'DV?�����l�	c���fɶ�>V���w�mC\H]|zl%��aʙ�5�%��uqP7� ��z�����g���0�k6��Y����4����E��A��4��	l�����u⤉�) a0����B
��.�[{#P�Eo�
([&A]�Ą��	���Eer���$77O6����w˄�ƫ�fz��>�fNs� � 0� �0@B7>$6��<�@���L,.�t�H��F����_���l*_�/�^}M������!Cu�2�z��%+�|RUfy� ���7�<Dbɸ�k$=}��]|�|�KKgX����)��6�-�X�����mX�^���=�-�DסkN���oZ`8���W�c=��3�}����m	%���l��)g��*|���xD"=�i�k.�'�F��;w�a#��c �`XMz:�<�]Na3�į����o�Ǆj\V�"�g����"P�b3
�l �gn?@g2���ڥ�2�����F�#�f�Q�oܸAΘ2Y�3 `�.����k*��@'�S�ZPP,=}��t6b����F�=�;jҤ�D=���f�V��}r�++�c����᰸<.����Bm��}��.|.\t��s�=�ﯬ}UmC�4g���~@U���*��{�J����C9gڹ�	K_����������6\���.IgP���S��ʗĝW)�P�DRnI��L���uIq^���=b��U_{��;~����
�y���_���k�g%l~�3�	��EE*Z�����n;&!�Ȓk��`��e�4��a�@��A}�1��,X,�9sgɬ93�ȥ�'���+�b���D],�� s`F��T� ���6 adZO�n��O ���7���3�N��<T��XU�0��xLب�\AZ���X�]��q&�9.����&���9I� 8 : ���š�Ə��΋��Y�@�?�,��[���P�H繐T�� �E��;��h>CD��8 88%��z��$��y�՗�����v��h����(׊�]wO��y�y�N��g����׼)O>�l�sX�y���)���B�����W*"n9|͢Yw���o�Rb=�l����~���G[r �F�]�;͌g�-�)���z%�I��C2��X��r�$���}�'b��Rk��%��&]<4ꢵ�U�#=2r�p���d̨qj���� 	�t9�z�jA� .��D������!MöF-����č��ơ���ͷt� �%<�ʪ!��.�Gl[H�    IDAT�����MF� u����Z���n�H*�4�l�p���P�Vq�iދ�B�qM6)?��r`��>��{��F��Ǧ�9�����x��b?� G@���s%F7P�\<^����/��a`'�#��l���<p�_t�o�q�\y�b�oJ�Y���}�E�"���O����d��e��eoM�Է�K��^��Ej?k��C�Cq�#"�͇�_8�Οܲh�)��t����b͋{�4e��xb����h3��Q�ϧ��X_��q�][2N:m�\�h�47T��m[�edoW���wTB�sLYRK[�tt�K,n6y�U�*���CE5�����W���'5�B�m
b]^}�H�_��J�TJ	~yyf�6͵w�Ϩ+N>�&�ŒI�7n�p�$�F�L> j tU�lI���SA4�5�w�<V/*T-/��{U���p^�h%������>K$��u9\�
����?��I����P�����U��	m�g�c���x�\uՕ*�l6�z�{���7� �}f��|����P�j�_���r��C�<�}�N����b鏚��8Ln��b��?r�%��������zy�C+V��Sݜ��~��"aq�l&IOj�s�]�ݔ]^��뒮�c2m�D�;�lii<"�jk�s�=*�Sb�= ���7�	�_����0Q�NDʉ!Y�m�W׾�j��4b����t�p�yPB�H�W9q'@�jD ,>�`�'L����:)K;j��OS7�bT�J��kjTHC�� ��B�`/r���y� :D4�r�Г����But ��ye��.�=�ZV�|F�N�BP�ĵ��	�}ҁ';=�/E��}qydŪ�ZiCWū��Rn����`&<�n�X����2*Ə'w�s��r��g��OV���%9�c�!�����W�}��X,Z��P������.�q��z����W�ya��c�1g@����]5�5�p*MƖ�K�m�d4"�xJ�%�=���(�'��E�Jw�qٷ{�><�m<&bs����Z0b��x�V/s"I!%���P�l�E�	�D��(��5��;�g3�@+4@Kj6� ���b�ϛ�F�
����I�iՐ���'(���%@CM��>t�I��j%:4Ж��qX�oX/@H��{@�����>~�L�	ܿU�E|kժU�w����a�"��G�1�(Ɉ��U�B9����������~_C:H�H<�=>�l��[�A'Y�,u���Ī5����Q�RZ5Z�	�=�$6�����Q��s��ў��m8�d��;�XO.q�cϾ�fס�܈ݧ�����,�Τx<���#a����>q�D�{Z���I�_0C��y�D�:���!Md9rT�Ѹ��sL���S���ր��ף�b1��	F+F ��ުq ��JD����L���z,��\$��T��1S ��.Qu�K��Y�+)3��h�ҟ'��$`�Ѻ�oHn��5$�{0��L�AYCg�*�I7���I���ܗ]AJ��J1�҉�� h��Ͻ^�>1*�x��D,)��'�-���?��.��] K��VG��u�䝷7�;�}�3�n��6�����w�w��Wٱ�F*�M�a�	�ʎ�{��Ϫf�n�L�[�	I�t��.�x��z�%o�Rb-��Y-q͞��*�h�ʰGR:�EIu .�ww*&���A������}NIFz����̜6E.�+Ǜ���i\}�:��Rj�kh�S���4 
� �asi����5�B\	�X��fD�Y��B��d�s�DD@�D��b���63-É���Tĵ�7���Z��I k���˪_��J9��9 �������Pz��Bb�q-��F��Pf �
m�2V�*�&���l4�Ζ��V�`������r��]{��� ���խS-����5r������@�����_�M}.���P�I�d�`~�8=9x�*ps�h�s�緻9��v�%�YW{ݢ��������za��漸� �_lɄ�I0�$����|�TL;�66?7;G�a�DL�?�p��9y�\|�ij�{�J�c�,0�j���tjŪ��^é�C�DZ0�6�`�7�d���Qj�U�50�2P[,8ҭƬ�I�l<Hy�G��� �8(�!���ݥm {Lal6�-/?WZ����_K)C�!�;�����&ث��sm6�<���W�O}�DVU�-�F
 ��g����u�vN��{B:!���ە���֪���Wd���d��g�-��)�ǌ��ol�ǖ�������W��$;�B��,�-(�]�9ђXXY�f�r�x�qIt��^�p�w��Z�ꕙ_���?X7�U��hX�I����zl���v5�����*�x�\�E{�O�	��͒��h�XX;�y\&}A�&K2a���W\y�2Nu�oc���N�."���	q�q�� N=j��e>��)��hHQrp��0z�0�9�c��؅ �HTS��J�ˎ��(�M��~�Cage~-�gY���w
'�3�0�6�����p��OLC1.�O�����a��r�`��[�h�|�����%}��:�q�]����i��)gM�o�C*��3�o��V>'j[d�03����EU`a� ����{�A�n��̞0����n��n޹��۝�`�/z��W���U�*DbY����C�8ER1XtF�љ���[)%��H,�#�!�t��K_o�L;{�̝}�J���>�V<�}9}~��/m&�
�����J��H���k����릱�D�X�7l<-�_�D^��G#N;��X[_��:�@t�wj�ic�Y�l�Ƌ
M���n7�N� ,�ʱ`�֒�C����	��,�aAU��˖~�^K)�,*6
P�����V���U�6��h9Dʍ�����j�~�m�̘9Wn��{�	ɪ��˪g_�#�M�/�J��3ck���bP�Rc�7��P��������j����n��|3�V�~��V>�җ�0�}�P�H,Kf+�X�M|N��"G���a3T�+&͍5RZ�+K�[,�F��c�u�a��RG�&��s����Q9l��z�n����`U2א&���f�7"Qo������a��c{!8yxzx�4��R���+�H����#}�I�sF���稤��s0�&a`�?ܫS?|X[4�R��p�)��(5�il�mFc�!� ۡr��Zp��`�o���������O����,]�T���-W_�Dn��M9d�3�Ȫ5/K�|Y����;��"�8(����2%�r��l:;����mW���%���p��so���Kן�x���~h�/��__l����W�d3fΙ�@+az�lI�S�,&����mw+����M��4�.�gL�k��ؽ�0K9�H��� ��7l&B�H�Έ��t���93��r�������rE���!��6c���2�T��I�.2:���D�1H%����W�54�.���d�^#�P!Q4=��k*�`�СU��A���mmQ:2�R�5�^�	�P�	���5LZT&���>���5m���ET��fLY��5u�+�����v��������)G�{�_�^�(MaqQq�Hjڮ��L�ZZ���Q)J#p�JT��i"n��a����qD%���p�g���߹��;�N��)������g���L���J��u:�b�|.��wIO���r���K��E|
�a�C"c�{�M�V�r��SƁ�=��ب�و�#��/P�B ����D�谨���FH6�{�E��o	i�P͜��A���0q�O�~�sO�*&�Cr (��������Ś�cb^��cb
P��!�|�6��� �4�G�G1�e�_"n�՘x�n�>\-k_Y+���N�_r�r�e���fy�����E��u�$�_*�LI�exU�4��H;�d�.�<X���>"1q�7+_R�er�n��fy�Ci`WS�U�s�7k���>�����<p�Ĥt�*��.�h��ˉX������;-!'a��,bW�S��5vJn�-�H�,둂�l���Er��)��gr;�Ӭ�(�y�'캙�
�S�T$i��Ѫ�@$ �0�?g�1Y���%�L(� ҂M�� #uƐ���7ޡ��@2�X��gΗƒ�Y�3��(�5�	��Xh���2��A���� �N�L{�y)�%�����@���TS �ռ������J(o���J\c��r���Hհ������G����ݛ+���s�'�T*�Ӗ�ʒb��n���CR���>ʕ=I��Q`ٜN�����)�A�x�Q��o�₳o��[���?��/m�����^�}����|��TH��$��k��n���N���H@r0F�#�pO�$"bû���.{BR�>	�"�ԳΑ�����@uu4��\�
D�!�1ǆy1��=j@��!��e����ץ�k �*�1b�Έ�9�KQs������Pq���$����B��s4-���G�-��Dc��:3<i����G�~�\�kX��lR��-j��p�|�c�@����M��7;��	�C}f�Br�{I�\��Z9���R�
���rp�!�h����K�%�o�I�/�T"I����3y��g��3)��6�����H�a�!�L��R�O߲�r��N�s$��@gU��h�.��<-���ݦ#\�^�${�.�{���|�W����g=���/�=�TjsfI���!��L�%�(*��ƈ0���żQ�^�X&�/5]�>�no~v:���H6�M���/�%3fM��B|���?Z'��1q���Ն�H��p��I�z����յF��� Os#�
�A����1�L5�G���&��-�����] 	)B�A~g5� T�;�����v���4����D1@��c���۷ɡC�ڱ���UR���U[r;�*Q9x|g�{���ML{i�G�K�a'l���=Sn��67�4�m<.+�{Uּ���̘d�|bw�%I���6��v��#	))�סZ8:99��O7@�W��J<i�`,T�j&;qB��$���p�g�t��.;u��ߘ��cO�����L�`%����Բqu[JR)6 �j��� �\�HI*[2"�h��b�����O"�FND%���\�I�&��Ek�����6}�y>��a�FQ}@�ZvZ[������6��a'�A��&�����S��\0����gS;	�D�����輑vx��5@m"���h�?o��!�*҆'��g�c�\@�{�(��^�%e����9ZA�TۡGi�tL^|a��z�i���o}[�̝'��|�������o,��"�$<b�Vv%�ɖ�X;����oV"e�@v�)��ln�l�ԛ���̫'?���W�T7���I9	RysX�c X�����
t*R>�Q2W���U���)���ɭ�=�������=���x��WaĨQ��aa�:ڕS������*'+����l�"�Ƅn�c�b{�e���xJ��C����!}�=��0��f֌�Ĕ������ !U���Ҍ	��ܢN A�B ��rl4��Dp1ǌ�> �E� ���2a�D=\D�Q�<Fvc}�l��Y�b��\r��r�e�ʸIS���S^^�Q��|EZz$�`�$>鏦�1��������TCYSu ���p@beg�h8:6"� ��8���"�rBY*� �Uκ�S:�׽1�/?�Y���P K�x$V2�	˶bQ#H-f��6�N���!�A���ۑ���6IƠ��HNЧ���5��ڡ������gL/S&MZW�9����z�MU)y���gkgAKR լ&�4���d��T��C��Qa�=�j��@-RH�a� ������K��S#�H15���<���ڌ�a�d. C26+L�\k�|���"���yc������u0�lI�;F!�<��k�a�G�sw�tv�O~�D�.�Q�M��!C8�b�(�T��HD|42).��v���	�bȦ���GU"� �qK ����U��|�mߠ
��zuOuS�wqzT(��- �����R�f�*��";`?�F"�vQ�*�� �)�A';%�IF�\v��=��m�/w�?G�	6�C���A�:HƎ*S�L[<)��[+����54Hck�3�@C�p�
�B$��	H�����Ԟ쀂��RC�B�	��!�^ka@�D9�Hk�!�s
<��|j�+m��th!��;T���E��u�<j���~E���U�k��ٯ�����BW
L���%�ׯ��v�������p��O9�F�A*"`Z0@��N��xL�ɨT�j�`�줁EKPKf+��:v傳�X+׽1顿?�v���rX)�I<�`ـ?�o�`��E�3ŋ�O&b�t���r�m�HŤ0/d����R\�/Y0"�ڕ�z�Գ�H]����f����	��?לWaaPrBn���*0ǌ)ϟ'١���z����F��<��0$�u�	��6��J6��PfL��k��kU�	c�C�gޯR'��3-�jN/j��l�����=����S*�QozI���d�N�KG{�|��]y��u�e�VT9D���69k�y�	����e)lݽWvTWK~q�$SH͐��̨N�?��H�0p��ƛK�{M�a���ⴥ��|kh��	���:`Q�i�_u�Y����o`7X�R��cz9���8R,4�2j�fg�1��D56��|L\v�e���&	�2��T쩨�#�2j�P�()Բ#��'CF��϶�_�(��G�
J�?�&�;׊ʰ��R�������UCd�Գd��J���Vban�ˌ ����H�S��ڱl:i"��@���K�-���#��<�tT�2�0q��Dy�86�0Xt�����P���̂|Uo�.Qu���:����KOg�Nz}���������O��.gO�.�8S-���7��/�ǎK��_N��<�l���@dI,�����T��Tާ��Rn��<�F�:���PU!��һ���++�+T��i����W�x�Sn��w������ޜ�ГO��{�q���x?�T���J*I� "�*��48
��&�e#�{2&��6;|�\&�D������|�c��T�²*5<��`�x���顆�@	O�{�$�҉�#����A�ԫ쏴ɘ�C5-O�jж��-Z�p�p�v~Ab`�0��0Ae�C�+[�i�r�a�(5�N����K2�F�E�K�\��yp� 2�>��J��ɪ�A���Oqi�aY�-1*�_��;��#^�sΓ1c'��W��.on�H֬{K��4�?�H|�\�%ą���1B6j��CZ#L�Φ�bL�8Rqq����(GQѺ��X_H�NS�	(w�*�Ƣst����ۛ.�y�-����oH�}o�_[�n���!b��gh�DhQ� Ko�N! �8�f�&�j��HF'%���?r�,Zx���*���-YA��ؤ�;,��|[6��Yz�6�-,v�_z�a�~c�;1IE�$��%p�s�YRQ6HJ
s�	����a:ǂ��*���=;�T�;���--�?��׬�l��h|C�0>	���key�C�]�	ɿ��b�[������ei���!UR5�R���n<39ɤklԁ�n٢�r����7A�k��i���c�·��g�wʗ��J�(xN���|/�k
�Ӂk4��ݦ�8Mi�M�8�G��V��#�g�_ʊ���	,�78 ,_(�|NM
e�(���H[��3'��_?���#Oּ����Z�nۮ��vg���`a��^���O�I���`&�`~2R+.NIH��ޮV��vȠ�|�}��2u�$q:D����O?�w?�"��S�9E"i�ݮ+��hQ��&��$H$���_�z;���/����&LT����&.4j�p<�R_�A��;�����9��x%t@���D���,��V����7r�h-ٯ�����b���p:�"���v�]{��A�u�t����O��=�KJ+$��KM]�lݹ[>���r�Ai˟��铄zz.� *�JHc�#��=}�R�`K�_R��%���@�e�d�W���h���
� )� ���T_[��3&�����[wBİeˆ    IDAT����^~g��{�{lݎ}�#�l�U$S��M`ɥ�YC���*y� _�V�yY~��j���j���P�G����S������H<�ӗ��qMz���MX��dB7��E_w����T1ӵ�qhh&���&̔X����Ə3P�UR�'��rhX�f��=���g���֧h:	��II�(ǞC�0^�O��(���,�uoO��V��C�k[%ʰ �Y�x�]�<������ʓJ8��y���DisI�Fx.�V��Y�Yz��y͡'D�Pi Z�F@L���d@��E���X��xJ����:x�H,�ǩ��ݐ�kkY8}�m���kO	��7�3����X��H�P$����&5����=eT�,�d[5�RތZ�+�\�&I�=Ӣ���Nm�&v������giu.R
Y���@�nI_$�iZ
m��X�ˢ�^��ߜ�u��,�0~�L9}���1��<!�p&U 6S4�3�V��qd��v���S���������>q��n�*�tTKO��낉��𑣍���&@[�9Z/ﾷY����;��
J����'_P����	^�`���0v��:Y6�gx�x�L�¼R" K� ���y/T������X�XRB�yy�Z`���?c����ђu6��4�3Q�~�c���J�".���4�H@��q�sBH�ؓ&1���)I�5�CP.��8�bT���ƻ���	
�fw�E���ѨƈB�^I�H�4�����%ĆS���aS��Z,�AR�HX��>-���� .)*�!�+e��Q:gO�?.�dy=:
�~Gw��tuIg��E-��so�{���>���f�$��qh$���Pţ���2�oϾCr��N�Z�x{�4�v�ǟD���aX�˫�.�$Q��X¦ײ���s�9��׏�N�n�a�a�-�
�����"�{4&���F���,$��p4��B��-LX�0�s����o��膵��Y7p�*LK,V4�VU�kiĪ�Z�J		W��Ї&��T#9�nm:�Æ �_�;$�c�T��C�p�&	��s"��ax:l�$��Hh�Kg���oӾX��p��$��٦��=��p?ܬ�E���KQn@
򲥼�L�����h{"�)��*qQ��g�{l��9]�C��@�V�HT	v���#����)��;Tݹ\��T�(u�CI����1�
������Hݘ���������ߕ!(�BR�L {at�J�	�B�qF#R�����]�*$	m�{%���b�a6Xƻߝ�xwKۼs'�>�����ŋMR5���?�~��Q~`���umU�Q&{e�*Ԡ{:@��(���s����IXF�%��%���	 ���D��a���}�C���Ρ��$,�DZjٓbw.S+�Jz�����v� �Nq��VYH$�pz���\��X��e֜v@��_\��C_
#��
�A%s�<��E��Qǵ�I%/�$�jw���ZW�T�jT<a�$�n0�!-�q�tk�A�t��f5��%^�!6ޠ�+�5���
�tĀ&I��P��Jqt��b0����G��<��v����fӖV�Mb���O�s�䊗gϞ�Z`�Y��������]�ǆ�7����E�2ExP<�#V����J~���jԛx�1���Ŝ�c3�9�0�|$$�K�c�$����4��6�8�nm�_+��cN;� HpֵYLT���ŋ�xIRa�r�ʔ4wk$��'Jʌ�nrq*�sڞ�sМ*�m̺�k��P��]&���PV�H���kݬ��@���FH��>��8Y� k���fTaTJ����0�b���e�*�؈�Q`�+�=�P�/WJ�Ms��������q��w��zy�������n�y���������x�e�7T����j;q��+}��x����$5i�l g����H���06�FKIT�d� n�y`8`� !�	�z���ď�� ��O&����Mɀʁ����N�O�)d�I�E���%�F�X�R�A�j�֊g�5���g$�@��l"���� �Ҕ����@X�_l� 7!�XXJ
Xx�:�� _�,9z����X��Z$�+%��Ǝ9g��ιæ��x�)���������vlޯ�Oܜ�4���dK�I�d]̴�����\�g��-��-�3mc�.�F�M�J-���CJ%�j-7����^	G�����-8鑸C9�Mg��n�5r�Qit�J5�S7�� ���YUNZ��1H�k�]:�k(<F�'���J��iڶ���y]���en�T�*�	P�z[� Z��8��R�ﳮ���L�
��EJ+7?OG3���p<9`��Ċv5t̞:���'��`��=�d���;U�{�S�w���&�&�n�8�,*�M��9��/=�i�nk�s��ǁc�ڌ0dQ��`��>�G��� ���Ӧ�f�^7+����[m���4��8Z��]}a&ZR�{�}N'Ϲ'(;ܫ234�n6�����l��8��#i�%�d�9Z��E��em*��5�t}@�{@�q���e�κ�~.C���Oڋ�{�*�Ӛ�$� �pi/$%`5G�X4�Qj�l�>+��t�3u�.�:��ٳg�Ҫ���q����<�tö=��)H Kl	l���k��ƫ VZm������W��c� �Y4����@��:3� 
L	zC��.+͗��|����p�C�ص_�#)�/�����ġ�:\��r&N�ٌ
�X�RnOH,�g���)�,Uh]G�Gz�^epچ�T�Z!+H�!��i�c���� ��h��,�e�uNH���T�N?3 <���cL��p���v��V$n�XN�^IU�������#���:s�?�7s���Ӧ�-���`k�����ﮙu���;4�U��a!�d`Y�&X�����<�e��V0'7}�-ᗄQ���Y^�$���S�k���*tқ�X����ʕC�M���Hg8)��R-�A�
'�h��8
��԰��d:��8+�c�>��=2X�z��*���f#͡���L�F�$�J���e~F�e8�6j��5�܉ ��߫�F�cE�`H"f�e�hm��c
,z�Z�,::ƺ��O��N��|Ѣ)��}��Z�iK��=�~۞��X �����X_U�'$��_�<=��Y`�v�?]+<��?G �R)�b����T�#�A��Sa����K_Aa�T�#%��˳�l��oo���QK�%�kU&����N��m�rj'$�ٴn�u,pd�[�O�$`��Ƴ@�A�W�w��9�j����!�fX$'K7#MӇ7FmJiQ� ��
�X^Hs�}�ѯ K#*�&������a�����K�͛����Bb��??�~���	x��,����i�[�2nh�*47oq�,`e�� Cb���>MV�#`�(��:$��%ўV)���{%E7g���Sϝ.E�U2z��ާ;�7���-m״�]�*-!�2��H��6è&#=,�� e�8m@Y6��ϧm5+��ß�j�~W�0NHn���u��4�~�Eg큱���r@j�.�W*&e�Fbx�yy���H,"��VJ;1��>;�0<}���qވ'Ϟ�sJ`����b_��B�w��$�^c�$�mc����O����x���n� ��>y)!,�a��-}�-�w��������4����#��=Gf�>_��e��Ȼ���o~�'�<J|�EO��'�f#��!��#Q��˺7+����	�kTޠ�i�Nd�/��N���zH���ȹU�c�W�`)�4|�e��0�9i՘�v��i��`4��V�i�Ϫ(��5,[�=��ePY���&i낹=�W�X�X�lz7��u艆*wO�4�?.;���,8��k��Χ�J~�����}o�$m���
��gz���2is��� K��j�m��q�D����{��j�h_�L3D��
dϮ��颴>'�@Z��d���ZO����KQ�0oH�)���p��^"l�r;5Uc���v����,j��
Vф%��A�y���+��MK��ל)���7a	#�1έ�<Y"Y��k�:[�O��N����ơ��#�Wme�G�5ȂJ�_�J�x�A��x���q�5��%%��a�}�xf2~�M�=�i��3c���p*`��ɞ���{����N�6F���,`Y�0X�O��2A�I/��{5�l+�����qm����x�ָ���C�e�E�1��ڤE��=�$D�[{���M��?"�U#�ʕF��͙E%�kW.<����t��n~:�)��g�q��S:��j:��s�#roI�L���T�Xq�L�Y��J�p�%��5����e���I� d�O2����-���<��Spp��|��j��U��n�tv((>76VCt�!?�p�G_p��~���������7l�Us�n��ɑwn"�N]�4ܕ��5�@�/,;D�����n�AĔ����,�A�\0�<���K����<ٵ{����k��%��\��|��k�7FA��9���m��V�]h�U2U�	ivB
���դ&�a�g4]Z, 3<`�~"nek��L#Y��Mk�Nج&�kI�5�҃����Y����0e Va^��cQ���f˾C����/�E�*��T��TNVh Xg�����)��~��;N	�_����>�u�l���nH�/�րWH r��^i��|X��l)u�3
]�b��g!�� ����&�}Ar�.��0��#������%KI +�Ԫ$RN-Ԁn���2�{*�ԡ3��7`0)�����V�LG�Yuz��[[tc��B/��/5����L՗)�4�^S�{վc�2u�i�4�#��﷒�i/�r�bKhRB��
Zcu������^e7p�Ҋr혽��!	�:H�E�/��y��t�$��"����͜���g���M���%�;۶���wO�۲��4�+�r��X1���HH5��	1"@w2��p$���j궧m��t�>�'���`��ne�vv�*g]�U�$ÝJ�-�~
�`�\a��*�p�kY���� �ʒ���*��4�g��-�1�Dg�
��$p�h1a�L1�����L$ӓ����	ђP��o <Y���QKMX'"�ֆ�>1�(]�Bm�ϭ��}���"��64J_$�R��X��yi^��zw�L]~�����p��~-�>��@�/���u��>��6�Bw[�Bt�DbQ���#3���0<)f2 ��� ׀��6�������62+�M��.lQ�Qe3!*�	�i�&Vx}�fz�f�+*���kݠ�z�lh��J$T:�	�d�.k�J��47��x!��P�����z���S�3ߣ��p)�ՠ��ā(��X���,��!�xx�˲� ���}]H��7XG�̎B'�k��@VHB��Ƥ�x��۠&�����=;d⋝-rڈ��.�<����h�Z`}���Яx`ݧ;����x�~q���@W���Xփ��eeJ,XV�� �ƢФ��q�ƙ��v-��oC��~&C$�Q��OAa��P�6��_:V-���o�������+K�D᮳ѨML�t�Ԓ"H��\,6��g��s�t�)ڗs_���e���f:�D�Q����ϣ�X
��\��R�R�Z1���&�ó�d6�D�|�;��k&�13\����;bT����ǵ���ƖV��̂��I��pk�LY��������ןo����*ܵ+x�������g���U��،)x��q��m�<1'_����i���S��:atZ���ܖޘes��m��Ӣ�t$�������1�)�k�>y�#�P����b�dI,�%&n�CK��G�p$&޼<inm� sj"�r9���C�JJ��p��2��)��d���,�k�C���P�#�>���ԑ/wHrr$���hK�t)�a�&�~���o<V��3��^ ���y�eb�Wg�H��wMKi��ܭ&�-��i�P��.��]����%��TZ�:���2-���rr� +��,G>8�a��u��Ư֖-[�?��ɵ�l�������I��hRɜ���qhѯ +3�jI$X�vL��{2O���I����5MX����5����$�ڌ� �X.��GR��A���%��D!J͘�Ȗ�
�����/!�W������8���3P)�^gwODv���6��4
�	#�nI&�O$eP�H�%���JT4���a`���A\�tXR�"$r�OG���1���+PH�����',�ή^����D U:���S`MQ����C{J`m�\���C���'_��.��� �C�'Ң��?Q`Y^��dbAK%3N�?��'�ȓ��+�9I�Y�8��j�+K����~=�
��]"�.�R���������e�=~��s��g�a�H�IQ]Ą� QQ0�낺���	E$�$�$�d�ɝs�ﻷ���u���w���������ߺ�}o8�������c�	QL|�I4),��bç_���O��h2��:�AD�[��H��Bvnܞ*,]�7���G��[`���Xthz�`�N��)��ǥ�ݫ{�P0�9s�b��E(��Ar�ֲ�+�^�O54&�#KϞj�G=���Z���z������� U�	2N����$yc���*���7�����<!d�@l3	vV���o_ѩ��\{����ӫON��yב+CH��hcjmͰ�^��<�(�6�>_Ȱ.v��ըg��83��=���2�Vc�B~J�)��Ch�9��C�D�^�s\F��C�FEUH�2�*�'�0� ��D��5�o�k�}̞YT�=�\٥��-F�BA�0��	oL~�7l���`�=�D�Y��� �6*���<���3��$2� )����X�j#ܢ1Q/��ON�H���h�|Qsm��\�c��"r�����{��p�IG-���ӿs�C���*��3}jɖ��FE���������f��%h� ����
�<�w���U�V�^y��[~:�;�8a$p>�ՙ�eX<
㮷�P�"������x��x��d�9�1BT���
�-��Uaܽc��RU�>-5Sߝ�E�ײ��X����wy)�l	X�t=^��	,v:������hP���;��i���aA}���N4�� U<��k(��@�	��B�Z�TMlW	R�S��c���	|��gpU�����3�7�d#�>��1	507e�*>�c,MF��v5��sqY�;$'����j�c��9�A����p�x���;yK�!y/�K�Bj��L
B(�`U)Z7�z�Gۂ'۰��r���G�
�-N6,��#+SqMy4K�PP� ��Vu���_{�_W�k^S3&�P����2M�PvE,z1V"}�P����V,GϞ�p��	�yɉ�}x�ŧѨ~>�o�Z������Gs��~���ؾ5�+��{�x,lVļ������<��8ӿ^��KV��vI�KeX��LF��J4̕s����^��#G@����o���D�9}8ڋ���:��i�l����P����<�Z�P���-�4d�h"�7.�0�F�Ԡ����Ad�cY�����l�9�G�:�]4�RE�=h���{���Gm�Z��T�暇B�t5�'�"N)&�����f��e��x�8�y�o<�ʰT�95[�����ʨ���F��u�9_��W�Fzɦ�´��o��O�9u���5W�����0��/�C4�e$۝�f�z���[�)�p�BL���ᵧ�G�zu�xÏ���{\���<.��,�;HP3��(ч�pUc�Ax�u8r�8y�E�ui���N��$TAg*�}�Vu�G�iQ��h���:���٪A���Ω��;���Y�f)��!꣪�̏7,_U)Zf~ңu��w�|m��BEQ�>�F�۲��5~�Ά�:D��S��%:d0Ԃ �a]�c�-�U��j�Qw�Y�څ<҅ja�\'��Փ,�	h�B'�����������o糸�����3Ͽ�-�6�c�x��G�ŧ_p]�ƿ���EK1i�L�@���	!����a�w�vZ�4&>}
��0�K_GT���8�H��f}zQ�����������k�����W_źv �KQF����    IDATՄ�T?lf��:�:[�շظ�١�4??F=�Et���sZU4W�d&TbR�}��A-�Gԉ2�k�c��hQ/�����~[ߓ4,��+���m��CB�f'�>�ǪaX��C�P2;�ڐva�4/�U�k�O ^@����6�u~}K��,��Ei�� (�AgD$�!z�a)�}�\��W���u���Oᇭ[��s��'e��}}z�F�˻b��e���y��X��;�b
>��s�C�A|a:���x���C���8t�$F��Y��	���=K��F�(/+�!���$���T�Lf�[��'Of:� �����C��/D�]��T�mmM�i3]4��5���gA�:W��}�꤀j}����U�$���2� �U=
��
4-H���%9�G����E�A#go�s�ƚ��1�H���E�$��!�XZ���Z'5���R͝C?��bGa͸�|oV�ވ#+��I"!�v�uc�����˱z�
|��G�5k����^{��;c�܇[n���^�EKW��O���[�/?~���l��eqF� (G�Rn�����D��9X�j5�9�=���6n������b������Æ�ߘ�ь���/��q��bFX21t�׆uT��v5�Vi+�j�ż��<��f��3�MTǇZ���K|쩅g����y5��и un�����r�ы�ͣfm�sb�fXDѣ}�p ��<O�jm�Xq�b�o#�ՑX�Z������_�����I��ڳb�M��E�0�B3�N\֩֬Z�������G���7.�r3��� ̜�B��z��pʇ�Y���G��[�8}ʋ�ǍG�(#93�r
�����O� *x���X��{�s�w��QF��3g|ƒn陙x���P�^!v�܇_x�h�^&�F��h�s�����4��R)�}U'L�f����l�H����PX�V�Yk�y����:X}�(tXP4��<�k�����a��d۞�AJ��Q��D�Hzq�"�T��Vê�>qê����@|-�\�����IM��y�۳%�
��s�c��Zt�Jp�mp��c�w�Ƥ)6l������&��u�ݸ���~��aɒux���as�ѢI�s7�~ر�?�.��sr1a�X�$�]���Ͻ�J���Y��B\���{-[^������)3P^FR*NDd"qSX��$���~g͖���5��?5����|ì�k�Z�R��\��Z><�@�G��V�UF�����Q~�M2��Mú�摳��>1H3,bi�,��#HL ~��ڰ4���}B�/�ݜcH5���y`@>�kh�h�?�����,��g(�
�`��#��ҮX�tfL��dko�5��	n�#G�$x���/�
�Vm¤�>eQ$�����������7�#(��W%o�9�w�/�A8l0艷ˏҒ����[q��Ws���K܀&�D��1b�z˶�GTTg�T��8y�֭��qd��c�g�P|Zs�.T�M�2�f$�F�ϲI�U�Fo.��&�"t�p�Ia��N-�'�����q��d���{,�|���U`�,�jYd�܆P�"ϯO�����Y�*��@�kT��j���;X38�Mk'�2�Q$�7���zt��u0u�t�%x��Ǒ_��l݆G}�y��9W������3f!���"E`��ѭu+���	��4`5�`�˕�wߟ���dKÙ
{�$R�Љ,%�8�aCn���f5�UU���FC��ą�������5�~�Y��i�i5HմME���N}ikU3#��5�Fj�x�<N3Y�����a�1IϞ8�|i2r:�B�z�s.m�{������<j�����)N�-NޡQR�������7���� �Ќ����1G���\j����d�4��{�x��`��vLL�T�6�L-�CIƑ��D�$;?|�C���H"=����)��F��Y�c�z�$I��
0��0a�[a4I8t�&<�d�&�*NI2�:b�t(-9�A�Ŭb��@|a?D���K&TT�`�%p׹ڀ�HS�G��8�M�R��jPdX57�;�gi�I������g�P����={,z�(p���l@�S��u�to�wϨ�#x�w��i��R�0Y���b)�$s%�}i&���������"�8�U]ܣ�T��u�zRs�i�,��V@�>���B��~$'������ݖ���D�"D(�0kQ��z�p�k��t ����hު�8o{W]�7��:��z.,[�
�*;l�ې����?�易����e�#BJ�3g� �a!�H�_]���٣�1}<2�v+TOǸWz��&٣1�J�i�^<c���0�[��-�)nZ�L���dXv�6���b4)L]|Y��1���p��G�5�FM�~�h�'B4Fv&!�f���B��>Brkf 8+񦓁ir�n��)��CO�ǫ����xq�j�	TK�J�^.I�;�ܤ%.S��E&�|��N塢r�ژ�vq�r�"�=��u6z(DzACzm4� m��z5��|�jv��&)��Ç�{�.#��㯰f�F�z�jO@�����dRZB�(���G�?�6('uL�:�Ƅ�;(NN�N���q���L�7�	����gg�)nl�HS��D�$���h�N� �*{��h�x�G�gCx�� ���@d3R����u�r��z��u]԰��e���sE-�vm�z;q�A�U��Q�dڌT����@#rL졊&i�~�K'#V8=u͉Α;LHUM����|�Y��s��m�H��z֨L�<�'�8[�{�ύ?8nsq
�8��^��;T�"�0%��j�������qX��fOGqq��D.��h@��d��ړR�rI��נ�TQ��Pѫ����ik��w�(��7��ݨ�Q�<�91!��y��Fb��Ľ]*��b�(b�Q�����r��U�!ݖX�	�`��������F=�lo��N�]��\��K[f�?��_~Ӱv�?5��B49������c2��3�bAb�[��E��\��*ɩ�"�dZPr�js����2��By�h�:��T�C�ݣy,u)���C9�Ҩ$5ާ85��t�R�q- �jG��i�!1��I>(ۣr����)�u�fi�>F���Ph�#���0@ΑB���0���h#�r�ȗբ����EG��H�c5�-��S����&U�'�z���67��h{i�d��h�A����3�x0�?������ne��H��eg�F�
I5�0۱�k��Q���a��i�;���U��YX���7�t�S�EerYIG���/j���m���S.�;�[�1tjn2F]�/�[��'����� �q�Qi��5���g���qAп���R5.��k���>Ӿ�qd,�����o�8����?�`BD��F;����?0��{��Xc���h<��/ט��%ь�����pTЬ��T�{,��	b�&�gj5��Kl��KN�3��-q�u��"�3҂�?1A�t�t���t�J��q���<�oV���&n�sr�N��)L"K��v�o��j�����d�T�3�-�����z>�I���yD3�t�t�G����C��sy�����rk�=�G�pY�V<�bO'��q/Y\_C+��|���q$��Vy��sK�|��d�s��2�c��d�gbģc�tq	�f3��Dĸ�����:'��٩�U�ִ<Z�����̨V��q�%��W�^�8^J��W�zT�"<��Q���}K�kW����u�����t4������Ln�'!!�M��JI�$�b�V��3�ׅ�Y	kz�ͻ{��~��Q����/o�}���`�"�Y��ZH��@a
`�Y S��S�b �>A�H:N�S�/A�ťe�<���F����
�h�,�M(W���q�jNE�Lg(]�R\�vE��yL.���/d
qU��:�>�JM]&�T�oqo��,�>�s�Eh��zl��k���šH"��\"a��|lP4�I� �si�g|��X>}y���;4RY�ԊO)]ذ���=:�]�G7�LF�#��%�,+iB�L0 ���R�*Ka6X&%%��as�PU^���r�����?�jbF{2�� �P�����j�
�ܨ����{�����5��E��-c����ѧ)+�Y�RR1��M(�j��ݮp�!���ѪY�i������
8z�$��*ƾ�q�LA�#z6.��U��{g���EUmD��w�ʒ�U�c5X�9N�H�O�V3,���g<�a�'��K�
Yg��j�*�6I�Ni�X3B�r��,�²�V���#B�]��T3V�>�����FI#�ijΜ	�@�C�ܦ�r�o�qiD�"�n�!��>�
�J�y�}���__�lՂ5�	�I���)��=V�w��g_���u[���EgaE6�����Ib��Մ@Ud'n��,w����a]{뽏o���UA=�MŔ�#$XLH�ZQVr��-�6D�+z��3�ߞ�JΠhGӱF��D���(:S������t����l�#JZ:q��|��E;��G�<q�k���y��ϲƨG�JT[���TM�ҦU�� 虒����\U���>���璸�v�|����
1�>���HHt0[���CD������R|��\�j�gU=�rXT3d�c��L�9�y㩅�p�ؤUyzv��%X�#^�8�:��u���|RL�/���O^|QL8�Sŕ�;)f~<�����#YH4¨��nF��A�l��6�6nؠ�5���{x������I�J$]F�pv�3쇁��a?:vj�NZ!#с����(I�D��Lx�F+��cb�{�Ɗ�T7�^�4�&~�Bd,��ś��s�:�aϥ҄G�c��@�2��1�`�jZ!�~�V�U�:��"��v��;D��2gG�F�CP9��LbB�J\��8�=^7¾ w �Di����1���l��GHh�x�jIaUo�#����j�<��'��Z2!-nu �jM��:H�
�S�N}]j'I� #�	1�G٩C�Lq��Qw�u˦<��{8{���c�����M�r�k�vg�	),������Ù_���2�d�q�b1��v�I� ���;:\�2��Q�~��a�k��������� �P4����dU��+ѼI#\է'�S���}��|\��̉�1U(���4�J!$�5 ��,�q���֮�7 Ö��L\9�j�V��k�{��[�GI�H+������q�U=��!DU�s�e�F5�*�Tω�p'�$����T�����L�iQѤ4�04�K�K*>�=^n�P���/�\�3���)Qh����7%4$CMt
��C�\�cE��G?m F����\	'�(����=�A� 3�	�E����KK�߮탮Z!��/*���F��DRu<DB���T�a�Za�%����i3�c��q��9�#��LBr���"�I5���(e�c������u��MX�a�� �,�F�:!�L�\�$�����Cǖ<ut���h�T$uU)�<)Hq��`F0�,V̛� ���lH��Fñ"7�S$ep�U����=PF�j�5hذh��3$���q�
8�|i��IK�֐��,�6��&#㽩=���3�fG�D���֠iLWU��\���ɱd�jA̝�i�p��3�M�P,�z*b�a��@21���F6h��ӈ?m�h��p�ϱU^f2��E�W��A7��~�`b8y�0K�)�)at�*��_��<ʒ��88?�1J*���;3��W�aLȄޜ���f�R̋���NM�F<q�ȵ7��_�a�$�L�_f��F$���(����F��+a��*�D�-��(P��5���1G���GPeׂ�R|39���X���tTЏDs���΍�	���K�*�MBĹ@���b�!�g	��ZH��b��P��鸩�'��s�0�W�&.+YHj�1�Ve��ܮ�,��f��~YYq�y�����u�#ƍ���yhD>�-�(S7���5�-|$��Ԧ�"�*\�G$�p\�Qf�Y�UD�hR��GǏe����^R�5uH,���;"S�p�j����lg��e�v��_���n$����Ê�r�9IҁvG==a̪�֭#��|�Ήި���V��,+B�E�>=��k���y��0Y��S�����ؼ���0���Ga���.^�U��dNDbJ2׍����Q���PO��Dur�b!fm����e�$�ĊM�ARU�)��D��j1��S�<�Fߙb:F�BFi�HǕ����t���ɃQ�^QZ��Űbš�P��0��P����E�G ��oa2�����1�A�LL8�s��悞����AR��ȣ��"a��S�N��I#b�*���Co���x-JNU�2�bvZ���W���B2+��jم��t$�6�/,��W�����ӓHC:o*��N�o�:��F.��a����k�M"�2X�p� Ѭ^؋T�	�ꅖ���+�b(Ug�x�2 �~��Q�����-I��;��>��箄7�g�"���Ԟ2EMo�]=	K��|�z\U��el�Dx=�jc���X�|��C��> �j�v
�{�|J4���*�Q�:B԰�!R��P�0%�u���` F�	N�X%g��n �a�:�d�%�PD=g� %Tz?	�i^�2M�(1�m&n�W�� ��H���;k�,<	D��ҦixDdJ	�E� #������x��	�ت)�N��plH�j��6�Y�T��gG��$}Gɒ�tVi���:����gp�'&&72u��7N���	c�u��+/C�=q��[^�:�ɞ��4'��M"n��Z4(́�_�JW�Q���3��{n���Ѩ:�M�;RMp�ʏwg-��7�2�`�'���0&G2q]>�S��BA��r�'h�Y�v���UI�N"c5xG�R�[�^����d�!�ޅܼl�����py�v�'��`&6��i~,�L�d�T�.-9wU�V3{j�P�6ǁ�G�#Ā��#��5y �Z�����A�|npWU�A���M�T��UE=2s���_���jJ�R"$%J�1�X�	&x+� E�x��'Q'=	����@8&3�ٸX3Ѡ�	,�b�ě��()��H̓N?���z����x�p�Fbz!#9�'>#A:ܱa�O?8�Z�W�5����[���]!,	IHJ�#����"�1�[��B��R��T���|ψ�����,��H*�_E�n �,�<|�3�,��#EH��KLE��C/�* �l2B O�.C8���d@���e��
/�È����ƉSE��{b
�4�0(��8����ѐ!�IN
sY(�J?<�E刉f�@�3AOr������I��<aʊO� ���ec���DVN.lv'��ڋk��ޒ�Ĕt�.�e
4�dHN�� %���4,-�7E�u��?����§�}���Cf݆�&����pa��dr$�}�D�����G�h^�X
<�
�j☗�,c"��j�P���('K��D�DoDR�J:�9��v�:L|{~9^gz��Qu?ө?ܶq�O�?��5��g��]��`�`4#%%r�c4�T����c��(>����53�Y|����7��c�Ͱ�s9�X8�|
�K]!���b�>\���\�ɣc��H�g#��v������Q7lF	�pK���W�SP�j_�:�Jo�%f{
'|�s;�Q	�]vR���nB"M������Q�^#��
���%U��d�Nx~j�F��`�Yp��!�$d���l���QP'��\�������I,\�����L�J
�:d�X����UE^��C����l6r-�k׮h׺	��8����v�59�����1q���ce�8�H0+�W� ?^|�d�$p�E��R_���e*��y+�U��F)�0BO�7��F0�AVN6M���o�?�J��&���H���O�n�8㞇���Q8l�s��_�����`tezF¾
؄(�R}/��/���c\"Uu�7�"�|�\z��*(�#�D�5�!��$%:�������R<A    IDAT
=�BJf$��f����%�	6f����:��٠0���?��0rs� � Yٹ8S��O����v��~�-i�*�r���$#%��C��	(r��N�ׇ=9?.âU�5$��3K���y�JQy��fn�ڬ:$%Y`�0Y-(���сw��=G���9S�jM�\�6J���I��"a1*�d����V���r�\}��نWޞ�򀄄�l��� ���� Rd%��A�_�ƍB�&��*;S]� .Q��U����,г� *��F��C�%zB�Y�pe��%�L�wP�5���)!�I5i_?k�#�Ͽh�>b��]�~���;Z��!)H3#?##�ݎʊ�\���j����Ү��NP��eb�H��­;�����!!-�E�C�wQǡ��Q��u���j�aB�{ˑd3!++C����>��[ɩY8Y�Ƣ��鑘����J�.��?C�`�B��233�Ч�d�����ȭ� �h����PqL�48�x��L&��:�:r DY@�F�eُ�yYHJR+�z�$������'q����IO\�2�VLb%�w�^v
rR�8q�g���s6lؐ�>��^�:[c��-X�y/��8C!�_�H!��2C��$a7\e�q��Wrq4	����xI�;���W)�IT�N�o��
9J�u�V���31���
�%�YP"d%I�;6�|��	�f��a=����6�#��-:�u1ȾJ�:ad�m@?��Aee%S&Ү��8U�)m7�-��AI(ã���JF3_�h�Z�]�	z[
0G�>(WU�䠛�ղ��@;0J
��w���
:r_ϙ�*o y����mc����������y�P���1���"���UW]�;߂��a����K��_u����}�qA�h��?�?�����Oe1�~:�o�˻w��ӧ�u�.Ȃ	!�PT�ŁC�t��Ʌ�Mz��:����QA�lX���O�=z4�6m�I_Ů=�0l�#�s�^~k&�IY��j�K�d�Y/�NF�f��(�Kø�#���|�Y���&q�2�^ D�|н�z kk� � G����f�
L��k>U���6Q� �)��� 㑧��Ӌ��><o��WB���d�`ѫc�&!��9)�]o΄<�~���%h�B�vS�
zӋ�5f��]�G^��;�3f}�-~�w
	iy0Z�R�F�(�W�~3"!�u�:���n�E
T�jѡ}�1���_�~zN>\A�T�a�xL�c��:L�a^*Ĩ{vm���F���x��'PTT��?|�ehݥn>
���;��3�~8�)�%����c���>ΨdQL�$���n�~���8S�39�v8	_X���`Qsj�����Cߞ�Ь�.6�]�#�ra�ر�M?���$|�x1F?�����ɟ�`K�՞�8~���p4 �B�݀�4d_�������ť���"8��4�P"��N��Foҳ��(3��j�#95�Δ���_a���p�t�L�83����R�v��|���_\԰FNxK6���B�Hc�`�$!�b��ꇙ�m�W���@�����jY�U�FR��p���"#�v�т��W�e�p�$��0��%��h����$�81Be�QV�9X������C�+{bǎx�ſC��H�)�;$�ة
�b:��)5��	�J*�J��c8~�g8�\wM�9
k׮�˯��͌�ݻB�9�e�/ض�0̖,$&��2���pX$[MjF�WСm3r;N�8��k6@��y؉�ŕ�}�9��Q��+q�W��]�i6���-���6m����y���p�T���gt�s=���Ĵ�!(��Q�yB9��¦�u���MK�?��������.E����/).���l1������$���7�@DeyNIM�39GN1�a��p��U:%F�*�/�H�	��5H����5���x��a�	�si�>B4��$�Qu��]۴宺��F(H]�ۡ�w�I�X��K��ԴL��{��O?a����{��-&R�⪼�"�nG�Q M���N��I6�0��Z^�����Ո]�va��]�%%Þ�ű�ƭ�Q���	V������TA�S��d��$9���UhѢ��ك�+W !%��4��k�G�9	΄<Κ(�LN������t4�f�-ѭs�)��c�����		�}�$~>v���ZK^���)���?�[�KЦI=���U������	�
��6@F���h�2,Z�:[*�Ss�r�<��r��B�!�$IV=���A	y���@�^]���l��	wP(Q� f�2
���SE����ث�J�/\��뷡�< oH�+���L�5!�Y�(��tꎷ������\<��Ћ�.�~bPtBoq��@"��(���	���@,�E�f�Ы{74lX�����! �@ U�uF�mNx�!�U�����X����V   {/8q)Pk��gt����>�L������d7"-��G� �����$H�#)Yy(�����*+�@ J3V����JuZ�.;���-��CVj"l&��*/���FE�;����;�x�Fk�K�Ф
��h�Y'���hBZ�VиQ]�%'0���LBq��vGq����T�����Lb��c����|#n��Z��n �U!�a�z��-��}�p�#/�De	i��b�?LMl"{-�!1(!$��H�造���NZ6o��W�D���z#�6�A�,�b��`5rkl��X�h%v�=��X���z�	)��=B~d%����>���w|sQ�5��W��d�?�$ `���.i0[u�
�b��Rg�����(�ָa�l�u�Nt
��O�����������q9V��
���"fJDDTU%4Qp�{���c�[��S\�uq�#�nF����˄�b����dxɁ�Ǳ}�Wx����(�ZN����<�NO@��u��N%�,����4
���w[vdOC�hM+����9I^:�-�^4���Fu�Ѵq=���q~9r{Ɔ-{�[��Ѧvu
,:�p9�N��K�gc��p��}9x��+J^hl��vb��X�~��4�2U�X�^���zO)8���
�@�+ѩ�x#*� tRi�ԯW��M#� �Ij��LI	>������YM����Q�Ęm`"���mϖ^�&����O��	w}{�둉,�~�7fC�5���Ov������N��Q�;��U䁤v��7�8��*���GY��.?\�²�t�z�4��Һq96���+@h�U3y˰O/ZvV:Ru:#A��?��r<p��I��a�MN�vƃqr�P�C�cO+�aX�
�0h�u�ݧ��_�E�Vpi��I����L�M�IaB8�նU�� "�"�:�����:�LN1屓E8r���}��@����D���8`Arf+O"�;���$t��
�4k̍���r��]X�~~�w&g.�2		�$�T���h��Hr�����H'�� բ=K��&�)��6Mިx6Z'���!"��p�`��J$�1��39q�Y��W�� �~�mô{���E�
~u�w+7�����#i�K�F�B�êl��`�!&:�Fn���Wm��hr:&��s��� #bn5r��+�<�W��O�poP7�Ԁ6Ү�	{y*���%BC���e� *� ���G��3"����O��#��9�bn�iw	:u�5k�a��_`����#�`Ic�*58���2��l3Tu�zOs�E S�%��Ne��,�@�,Y!��@�3{,�w��0�d�9M�C%pU�BEe1��:xU`3Z�� ��9a��'�Өs�܅��Åd>�8���Q<��Ϭ�a�@OO��f4�rOPO��(�����E��pb���$�cb��d��b1�f�	T�0�z�]�̻u���C�hͶwB�����T3V�gR
��,@��.�4�N�%�l���0M�Ќ��}��Kd^��^\҃*�ŇR�A	*_XzD���!�<4aR����i!U��{a��z�$廉/y\�(i�6��(�q���P%BAC�	0(Hf̉��6�����)k"z$��"��#���g�:�++�r��T��6��3'����&�Tx2t�ЩL`ћ!MT���| ���<��:Xf�	�Eup�ɣS/�	�5�cI<�x��h�/��h܀�=�>�ť`�R���O��	�D	ڣC����NFy/!G�ؖN$���YB�[��L뾶��C{�5�1����������)z>�
K�MVM���,ԉ[�3c��$��
����0��'��Qˆ!��60�����9��xk�周�-J<K�O$������A�f`z8$��_T���"�0Z<�Le��8F�[#��"�SFk��C$J�t6���P�*qB�JP��i�H�t,f�D���Mӱ����EYx�4ED=P��Ǿ�-�"�H��Dj!�>Ӄ�"1#\E�43`��	����3�&�5�������b�Q������u�֠a�֐��u>!	'�ܧB|��9z��f��\�&�3�D~�eoˆ�?>b����}OL�n����?�?�$�*ɟ�aiHKY �&u*�0h��Ӡ�<�̼�q�L'�G"�IZ�-��ş��S�"AK��v�vO:#Y��P����~������HIA'�`�� �iV�NG��H��^e����F��G6f�0�t��"&ze$j�H1&�=���#����h�ӆ�������@
�	9>C�)a�������c��3�P����qFCP�G�1��R4E{�n��o~�ٱ!1��g�3���V�ɘ��RgV[PL�MY�H=E�z�z�`�2,���O����w\|`����y��͋]A���@���ƌ�x���S�_�?�6�Ju��UQb��8�${ �k��K�,��Ƹ��Lj���u��N��O���6i�[�AP/��$D���-�{��3��P$��~6l�р�h�����Ltp� D%����9Se�%�D��9�T	HH-�Ř4&��F����JTF����I�H0�TL�	�Bs���� F�T�R=���x°3<L3��k5��5rZ{un@�gMF��P�֎��,�!9�1�J�'��}D
BjeF���0�߷��8�1C.��E�I��.Z���J:�@p��C��.�X$*�� yyF]��T�E'�ׄADAT�T跨<�J,*+1��Y�`M=M�����A�GeY6���&BRhA(�Tb�Ng0�F�^��ubEE�>��V�]4��X,a�a4&GBaQ�$I�ɂ��b&�����c1�� %3t�Q����7%��AD(�aO�~?�S�F�G��:�Eqa���*m�,��'�;�-�n��R�H`o�2Q�lzE�	��yAc����QAb�qj.G�/����j��X^�*���zc4�rL2�c�)��7(@�Eb��~^L��L�h\�%�?Z&�C�.Y�ߟy���BaG,�Ag�E�J�^uz�$Q��כ$�"I�l��%�)���Nug>ӣG��節~��'���G���,�1��3�"�bQ!�2 ����3�9��bL�	Q�u~uQA�����X�Vd��bQY�
Q�C� �1A�f�W2(�()6�5d1����g٘��BP���)*ʱ�����`0���R��M�:2W�H�MAg�%%,����P Ag0�}��$%��z��(>Q\�h��u�3�z�y]Q�)QY�ƢE���2:�_EwL�mr4�0�L�٤���c0$�&��>�N*e�hBVbaY�I:IW�Κ*a����ɒ^�b2�����p(����Ű[����/��gE�z�6���)zJI&�	�DA�J�HX�E���ڊa�3@J��3
 "IBD
��$(���(��H�bĒzoN���G�Rϧ�����k3?*���)���5D�k���_oC�#���y		�m۞��7Z�l���{��Qg�L��Q�$I���XZ�%2p������	e��4�� 
�2�t���fumע��w~�?����a͙3'm��M�VUU���c�뮻��Ts���]�j�i���,�p���L[��}�?���=���̸<��wj��?b�t�w�M�����6m��f�=ѨQ�j��?����|�_ް��ꫦ�/������G��[n�����.�o��߼e�Ċ�Ҏ�ٹs_z�񱵽�v�ԩ�y}��~�Q�F4Q�WQQ�勯��T�c�ԫ[�缼��[�l��V7��/���s�,��h��f��Uxn���X=��{��������/���������S�_+��xM�<�%����+�ӢE�#��ŏ?���t��f��K�����yw4m�|^m��g^��7���5�����P$���*t�m��p�����"�wqg��沵k�|u����º?�;r�e�;��kϞ=���V����sX�歫�~�8�2��9KEQlոqc���[�4i>����?���Z���/?_��nw�����4xȰjP��]����r՚/�%�+�����o��iӦ���~���b뼹_����.��ux�6������)}�eKcr�y��]�9y�6o�zMm��g^��7�-��՝�٧K}O�7�����!����������/�Z�fŬʲ��F�o|�-W���hϞ=��W/�B:w�4�M�N�6�~�)}횕�B�`�ƍ���f_޺i뽿���'\��7����gM�5kYyiY�`8��߿�ȡC��:���z/^��S'N85j�e�]w�hѢ��j�"�5�7}~_�n]�oӦÂZ�  ���+Wʈ5���;^�a�^��49X�������k��ԩS�.s��-|>��O�>�F��Am��O?�l���E�N�7n�y��^�977P��PF�`��K�~��]��նm�Z�{L]�d�ZY��d�mT�A�K.��Zd����ϸ�/oX�6t|8���`�mUUU��=�7�]�i3>�x�Y��Ŗ&M�����1��ׯ��}�c}�ݼU>��n�]���<�K�.�^�z�Y9'�����������w����'��*�v*++w���Ə��a����^˖��_RRbjԨ��{G��ִiS*Q�מ�=��6n��=�;u��S�Nsj�v�t߾}�KV��"�bAZF��zt�?ê�*�/����w�Z�������]�v�����Q��N��р�˗QQ^�kР������x�C�9W�^�����w��axǎ]j��ٳ'c��U?������z�Q���Z�������}��#�x��K++˕nݺMx���_��Mߛ9��U�W}�r����
��wϘ.��E��jՊ�>�7�]��#:w��am��Ν;�V�Z�U�I���ig�7jԥm�f�H��ߟq�_>ƢE7n��Ғ�>�5�~�e�x�Z��~x���+g�=�7���ޱ�v�#�U��}��5�}nO�v�;�ձK��k�`ɰ��\�E������Ӎ4�ڼy�jɶ���ϸ��°{p��GO�����C�=&����j����}���+V~J|�
�����u�ܹ�Y!��������mݮ�m]�\�um����+7�t�:y�9��/�ڢE����ϟy��a=��O�;uquv����Gz���.���s�u릓�����;ꮻڵm�V%��ŋ����[�nuS׮]�9�~�m6��S���oJ�:�s�3��׻�u�������	��w��||�T�mD ۪Y��x�'k��'�=l����'���ܼ�cGk�G
�G�1�\�r����n۶퍝:uZ^��yϞ��lL��


��6)��ma�����3���0��{������qI�K�zṧ��2y���o|��v�n^����tN�8a^�x��ϗۺu끗^zi�{��7��X�t���V7�0C�����k�����+��7^�����H̱~��������v�^�<u�7N�UT�NN��Kҽ  8IDAT��Nhݱc}��/2�E�m�z�mڴ��{���c��6��oϚ�`�K��^VA޺����������/���0�7'���}?=������5���^����5iʴ'�l\����rr�~=vL�V�Zŕ�~��6�aÆ=qú�{��3���+�nݚ�r�7k	��9vԹ����FZ��s����W�;Ӧ?�y���B� ck^z����j�H��|[6>\Qt�ٙG�=<�M禝+j{��/^L�U�m۶Cz��1���شsSΪ9sW:��y[6l�������o�~�G��[�����ᰡI�&�_yib������za�捏W�BVV��Qc�w�СCym�C���˗��}��Cz��Uk��j�֔����lw�L��XֶC��H�����y��ǚ����-\����h�ԤI���=�z��.��S^{c��M�*N������n޶�m�31B&,X�`�����ԩ�m={��#u,��Y��ٝ�dfdu�]����������k�֭�]%{=Ur����	������<�w#.i�jә��,V1Z�f��p�a�����kU*X�jUBeee����ddd<ݤI�ٵ���\�$�h�w��&Aw&$gLMO)ܙzm�Zf�Y��6�e��:��X3�T��ۂ�`A��Ѣ'6�_2�	��k�r�m���ff���;O�y�x�bhH����8Ä鶤3�I�t��4e࿨��ܹ�:eʔv��q�ѣG���myyy���uu��e��_�|�޽hP��K��5KǄ}�}�H(���d���r
�m�vN�~=������>�/kXO|�~�%�>����zz���tP,:���A�Ɉ��O�%�{��ޣ�%ek.���>�"�����g�DP"
�Q�"��wkX�5�%�����	=o�y��|��7����'lڴ�{$1�"��4�G�AR-k��ǌ�#\�^~9ѷy�åxX*�����F�E=d���/|�ɀ��v?���Ai��/kX7�̼á���� #��Q�Tt�D٤93��J��g�;�M�	�[��1�o�j�j��[,���2���J�V[,�@".TD|142&vK��C��Ϣc��g�[�p���Y�YL���`,#>)�F�\q�s�,Y2P�S\�(f]}�K���M
G���)�I�P��Y I12���a�7�\z��ֿyF����[���-E�ND���P���k��������/���/~�n��j��%�[z��']�ȫ5�ƃ�_}hC���� ���[^�X���f�;�O���~�Гs�/�U�lC�L%z�6���ρ<�5�)��$	�H$"�~���:��=z/\�0uΜ9�?��çE1��ؐ!C�2e��/����#��c�!9�ӿ��f���0�\Y�i�o���6w��D� ���������֔�G������_�c]3��׎���ЧQ�a[�5��_:|��Ϯ߿���;��ֺ�?�x�`m�}��u�����۝��]F��p�����B�{�Q�k��YydG?�A��p~uC�v#4�%
�_|�U+֭��K�M7���'�|������[o�0{����a�k׮����{���y�]��ڻ�Pď�����g�|����u��/N	I[�|�����'�']�3�77}☻gâC&_gCe/^}{��IW��,��6�㩞�N{ж嶂K���qK���K������ue:�-5h����ݜ�����`N��͜�Wo���_^�Օ��������>}����˖-��ѣǯ*�.4^}��Y��YYY����K���G
Wկf�L�5������F�$sd�/�	C�\��?͒Te7��y)ۻ?0�O���J�$��͏���C_����b����@�M���|댶��m��X�׉I	r�)�:?�O%{�����^��,����N}?������q�rw�� fv�hܶ�S=Gr��\2~�}k�`RQ�@��Xi�-z��rڴi}\��I����;���}�_�p����<c�ؽ>N�8o(�h��4��ر��������f&��i�E�r�����9`t���
]���.�Oީ�@FF4�����Z�۷/Oݼ�jz��O�Y[��eu=u�ض�m~9��|�����g�GBh$$_٤M����ʟ5gΜ��Ʈ;y�t�(��U�{���~�7�|�p뭷�������3f��z�5ל��m����=O�����<�DR"#�M/�{}��嗆�C�WZa��*ȭ�2at��Cβ���}���aї�;���=CD�����{���_�#�vM�l��II��h����5H[�/���M����"!p�?����/���-n{���Цi���w˽�\�@v�Х���cwϗ_ƽ��7+6��k��ѷo���⋧Ͽǐ!C��裏&ɲ,���k��/�|全�����S����X�N4����M����uϭÏ�\�/  إ��!���O2����/iXc�zq��%���E(့g�/]��j���v���o��}p�u+�-�	��I���>����nx����_�tߺӻ_/IT995��v��F�R�yۏ�~n����ǖm�4�T� U�DGs��)�<v������7�z+��~r�رcz��9g��%˖-s~��'�͜9���z���뮻��2e�'�V�r��K�N����ϧ���͒ur[�����ܹ��O޹r�,��L��2�L��a�fڣ��d�Zw}��;'<��2��/����X8�y߾}�N�t=����,ʬ�����Əv^�ɽ��)��&������3��<|���32q~�
����A�O�A�Uഏ��[�!j��0�:uڴݻw%��������t��?@�	tp,˟?�����޳gO:�f�����G�'H�r1���t9�?F����9XE�~��󟝅�'��^U̶]��`*��d�`�Ιg_+z��!�=�o��Y�������������':|R����W�d����L�;��r�s�O)o�0|b�� ��
T�q|�ˠ�)����y���Bw]P֑�����[�"s�޽q���?u��������hA\\܂��t�9��ܳj�ė�GR�>�(����t���٘�2�g�$���ĠB��e�W^ɻ����l�Ҷ��ؗ�9������>|�j!�ǿ����Wj�B&U<�d��������������9X~��(��U�S�t���NGm�F9z$�_�x���իf>|��翧��~A__���)SHZ�'5��߃'����w���)/�e�#*+]�O�D�B�]C:a���Q}��фE�0�6�&����h¢}�HFֈ�v�{ �ߧ5��    IEND�B`�PK   w�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   w�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   w�X�Ki  �     jsons/user_defined.json���n�6�_%е)�(��s�m`��9�@,H�J8���A�w_J�7�HT���ʦ�oF���z������Q[��Kj���i���ڪ���]�1���[��ZG���?N�}7��mk��l��\����j�mY=���㢱Ua��2;��ˋ�:�Y��6�ᖙ��v��k�9e�C
R�H�%@��A�J2q����֦�w͐���_��rǩH5�@+, �TaY��Z
���wŭ����&i���	�"h�2 ����3�2b�~�./������Q��o�z�UO�r�)BI�N��x�v^>vג�@�Ê�E�к�������*u�w7�u�=�I���R4aq�a»��Ua���M��Mպ��*m���u����9>��_��}�?N7� x. p��? ���wn���r�c^��|qCU��U��e�n1���,l�\����^��ϥ���
�����Q�����W,�*m�<�:={'���T�+æ*�[[ͪ�T3
	��A�)4@A�]�7����$�N&���.]�#��r��M����_>{�AϰT_�e[�(˘M� ��! ���Kg��N�.>��f���4�]������jgA�s[���\{�tL�AT�g�1S1���d�?�#(�A�k7惊1AW�˔c�G��_�cY��_a?t,*V�+⇎%��jE�б�pX鯘:֓�������~ꄢ` v��c'4�°���e�pwN�h,,D°4S\cm!��O4-���O�B���O4-��~�D��T᧎5���!T5�Q 5�S��Aտ����E��O4.H��O�.H���L��$���h^<�
}���Q��$T�`P"2�����3��I	����G��7����;C�~Wt]9��ܧ7��ٚ��]�xV��]��q�%��:�[�}��m�o���Qm�L�VΘ�z0� ��1W'��U]��G{u�ɠW�9{�p(2(�)`��:���FMe��y��w�,���)Ԁ`�b&�9��pvʔKL2;z�2a��@ Ҁ*��N�X"�q�p�������7h<�A�)��h�8��Üf$f��d�8C���`�ȇ��zMA�o��o�P��,�����7PK
   w�X��m  �L                  cirkitFile.jsonPK
   w�X�<1	}�  � /             �  images/02d8db12-ba28-4e49-8e56-db179b980a39.pngPK
   �u�X+���q6 X6 /             d� images/1f8ef630-8a1b-4a9b-bd39-2911f79a26d3.pngPK
   w�X�w3.  )  /             "� images/b3ba8064-1e10-4daf-8b84-7882f41f3c09.pngPK
   �u�X.D��N �M /             �  images/bb8b4d0b-321c-4695-852a-55709d7923fe.pngPK
   w�X$7h�!  �!  /             �N images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   w�XP��/�  ǽ  /             Aq images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   w�X�Ki  �               �# jsons/user_defined.jsonPK      �  1(   